// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:25:52 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Pl5sqKC/KttTNksbAFA/zSZU7iGE9fdsVD6JGzMdxKdifNpSjdqWgtj0sdr4AA7v
1f1gAs7oSN7oBlkjT6acmI/wkNbwoBdkklpyz8Q3S1XN2Kau1Mv1BrvPvahKY4ly
IoSSoVIy3deTnK882yaKrUs+oChfx8GCk3PHR1Cvpa4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27216)
NYprs2BIRza7wTmmKIT0xTpIFP9LQltmeDq9pmsqDtmP9qkDpirpAYZjOARdhVYu
Y7DnJWBFpQrVgsGRt8xIWzF8jkqIIUFO4P8/2yeH4ZdMGQdjdnbf0NC+VwRQkoyK
1E4CjqOdFKCSkRf2oTTJ9NacWvwfaE2IrX0rXjtrxzkbBANvTSlSt+PrdaE3cEu1
iJ9pLoabQag3jQRXN712JiQfLeEmdvsaiOfKUi7D6Uzv/HpucCZ8y9rQKJWLQLMh
gOZYCPxdvwTPnTCc0ArmIJ2rl48oBLKdfpOxyCjt+feb/rgIH3KrO2Ex04Hjudbv
nVQFN/KCND6nEEAfIdmUnVPv+Q1T8HWVWTJJyG+6ifvgbIVz3wgS9kWbCHiAwkj7
AFDTo89PncqfuqZUKeh8ReLfLcLAGkvk+ycGpCZ9ZrG9JqwIutm7WJHlg794skqf
6mqoqEQKClCDinF5Ha1fJenK/SBRA/J1BdZpuDZ64DOw58YUjkrDH4kdYbTUBCc6
ZeM9d8O0O7oGnVai/vL88F3/1nZj5tmL0jFh8UWY/YQwBGZb+9Ce+izEg7NQIoDI
VsXehvM7sHuUoh2C13qqKYkmXfb0OCf6Vs6TcfanEWNm14zqyV+W79aYBooF6bWx
fhnC/1/QjPpA7Boj//OFI/CRQQFlKc0V4skvv/e+Zt94bPBneqN6KNOkFMs0xt/J
qdDUZkn2qLccz4fzL2FmcWUWd4Fe2xj2fes6K3kBbKkVtxnSIOxTvl8F6Qu5ACMH
x9J6QGEiOd/hz7ryQw9eb2t4W8hpnuwNsLyUhdwoXDQzUFgAjhkXkKcxNk4gydo6
+iL2KiOgr0CQtCOeUZJYhlinJmf4qAjna+59aZDTi99f0TDmNfNVE8jO8Cj+Jt3u
7wW32XqVuS5dRygQhfXwv+S/MaTVnp9bYb++5LKbfnIJOWXx9Ulez7RDAle4VuL6
aSNaswpwI+fWHoWHdBjUiOuk9MOZpdxXn7MR0GK6QR/R0mmYHsWZuBhScj8tI2xo
tlfQiq8LfvTxYo/xQfGsPNSIWG1H4FfGpJkbzTXECLoJVDE48W65z89xiUJHJHS8
FHSoTk7BaFieECV9iIB0x5akZP85Ch8o/QAStILalFO04YgJWxGJCCPH/gnuRYD1
ka167T2K2DvUVnP9soR+7X8SacAblkleG2szMi+8W3SZy2XbTfgtOBWsjRr/E/8b
CYmJ85er9gIEOwUB4vZzZ3dRDLeXCsnRqRwpSynTgyCZ9G9zSFR59EzSrtbklxFm
QsqhY3jaBrLoV/wCQ+q3+pxv/Jq0CZC0LQxRlAnPSJmwZ9a/2MkATJ9/5hM56CaC
wHTzomDA2/cIW5o9uE/kq1SvTbSuUYP+6abqrCZ78FaU6jcXFo3rybgQg4iz1XKs
B1k0Zpm6tJA9ZCig/Za8YGLZzuR3kpMoC2mVf86NmKiAkYtto9pNNPmvQCF/BV4V
j4zqVAeja1chr2Tw5nrKQln9Js9ch1xREEcBA9mvlN1jzj4AYKwAQQvaxOHeB4RM
J8kd00APOkbkYl6VM8HuJk6IFuoWYFg9RBQjPcn11PAkWsXWxs0GrUa8JN1ks09K
Mcb8SFoG5VtOXRa6fPEOz9oTYVX53YjAyBmMi3jdDV0UOVoQT1vxyw+AnHEAg+hS
iJoLLvidc+EYAZZVJQE/FjPFxJQk3hp9KfSwjEDmXmLNGlw5p17uQXd6i6yO2Hyw
Ub29IV5AYpRoLNfhZ8sPTCOUno/BWitZbv/Xaz9cZuO8UmCRq2rvSHBREBF5Dttk
X0xt/R1CokMbffTpZ8GkRWAld8uH1vRm518cx7CGrq36/CdCLVkF1JScw1sVM/oo
4gWG5EeOni3Ax1bOnZwrMKp8gu39Ldx6BbcafFAXo/iniZRMWmOHg49oUr8QM/xE
BcNnbpdrp2bSPG+/NNIBMoR0d8JhDuIaRRsZgRHYI8PARET8cOS58yqqb/Dgb+HM
hFMFD9Ak+V5Gsflz0iIins5/7wZn5c/2zD3SbHJJgkIw6wAWl/t0KD/Vf8GbANzf
pDQDBVVyR4K4ypMSA/lS8KsKYaWXoxFRRqFILV7QAyTAakhuYYI+y8BV8wl1yTWK
5UhbdBd6r/al1EQow2c8roGslmR4hg8LLC4up2x17AQRFHf4RNSiEl7gS+jrORxx
93+b9/dFX2gGUecMmP1meucnA3SgTkBmSPLDOSAtkShHRxArQfL29M4+7rTQnEQS
ZXbQ5EkGu/rnmKXZyOxyzVwlyWG8hNA7aWu2JN9CmBPNdbOADTnEw9KwgEsbi2Nh
zwzIK5RVk7wqFHaevXa4gaq0IsZT9dMozjoZYpNVKm5JVfhyaXVKyVjpbQ9KZAfH
0HQZ7Nfr6MmEkvNMxFwFXw6xOLyMs/NCLGYljIJhIL1noiCKOwgyLXkPsGj6rxwM
3Zm4kQMemvbfd35ZYDrQo6xijYj/i37zLYfLGwXOsggkCE9GT3LsyCcbL5wJroCo
tzQ963NSVLfY9mqUzWCQrAoYsogQ0lvS0WgCLxps2tsdy9ed+OBxI6il4YHuiX9U
vMhW4Z+yKm/oYsfyLGz2pHj66se8qYrZWpWzrHXtu97JHemckyXsI7EY2tGxUw4P
nVLWXVzc0SY8w82Bu9A0x22sAxWg+1+IJjFEaeruKRIexFzCpbgbztdPGTAbHKw2
zudtkb9Kg3J/M6Bw1MEQPQP9l9Vsqi+rqO8zJiLBMpLHebKINYZgmI2NYrvfuHdq
/554AZ+Ou0rh3F3Bb4+aXfyI470Kw0WIKcum/hDYlsOHN0RdUIRjwjRAtJszel4x
oTVgFkPauwwh+JElgMMSCNS0M2mQvB+ylpWi4/aT48h0DMkj4hP/6rjGicHA1eJd
Qp2YWaGR2Xs6mQkUk5Bj62nnpiaq9M1j5yOVSrKKJUDnZehwf3eU0w6t2Vd4J077
NiMVKMFH383JhZ3g0npTiS40XeJwqiB5MIXgRIoxDDRTSfKVDO3jaBzIh1qHmoYc
+sXZhXv6OJroBamim4DMZUFrzi6yHs4QauHK1hvmBuPmzHe+1kHy3rvnO2Xvn7Fr
Jw5H8O+Vqn9H9+CKbQqr3xVvNKhHrADuMYwSAGVp2vgAN4IIBMXwGJ74rjZo4QxK
BjZGZeyB+JFv3iUKBpOnyXF/cqyAbdis9sojdWSdjG1mZhYb0JT57ObhRVk/wirQ
aJJKnVuWQPMBc6hUNDLP/s9/az5s4xAAYqeVp12KBWbx3YR0eddH5ELBeM/DN+9X
Ec6Uu7gUogMM0/AbbKn4WfjVKKms5pWAGmRMzgDe1Ou57/JEw5XBIyLQQUkotCef
k8w1Y2k0vMZIii4bqZfjs8Ox9FV/BPgHgvqNOwBqBVcdrEtumBgg60MOhK6V38a6
UlMINUkdLtRZKYUyBVbdmc/8psNUyuwc1p0d6kcwxBgzBznYjA+Qck0XQZJ3bgnX
RbYTxLi4LkNGKeUg7X0oJ0ashA/cqVa+c2/3LS1ELqAnad/xcqFjO+lZ7AxNKxzV
7kjGV6pUo4wEVZeHeACi1WPGbiwvykh+lBnNdhk7adcOhWH/cOCBEMws/C+eQGbG
Xu6HYU+2VNwF8D+HTw+morChfU+VYKqfI0cYW7fF2+DdpVCCuDtO87NAwG+UYUzX
aMKHL4Eq+BP+Hdfh7mca8MQnNUJ35s7lgtbRHiDRWgqnxRI7YY5mplm2p/kMHq4Q
eRtOoeXPbmT4DcscWxUFcS87bH/2nznTGqEAuAPLGvV7RDzNUsPkGo+FZmUtlFDz
zAWueuCPXHZ9mEk5FkDkwgihPl9evDDcDSu2h/8ocQPE9P2bMchEK0rbqX5ZFtEN
nBtW4R8PhnXor8C5x18mxu6v3Hz/5glXCwvNpjIFu/xHIZ/EJfDgCNWq4WZseFFq
G7JkIW69PiSQJKa2F8k/w5KJaWoIoYPcchAgidsck2nGIQZZWDAU0TT5mR9yejmn
Wspa6jIiHIZquVr6BEVpMFbdh2M/mY1oi5RwGJbL8rRa/v0wSzZMx9ogTEQX86Mt
yI1rBhq/Zx16seU0EqH/iZwG/vmtlwM3a/1cu+teiaP3+w5MR+7tCIluhd9OQgyt
wmX5j1ZbFvgI1KZ/O6NG/QOl78OUJ8HmrW9WracmiHs08J3IQGBTenZpnjVphb+e
v3GofMwxEmI/yWv245quobW3kNgCjdwxrDRaQo8gGrBV81RdGMUYf5KO9/4a624c
L20Ak6Qa0dXBIOf0B5pivU9OCID6f/UrzdJ+qjS2Kd7qlj8NeYq+HpKsLsvbCIMu
71yu3lImt4VC5hjKYDu3qnmt8Ov3IV5+VA/ziLFBZ/2av0iSYTBFpm747zfBcpFp
cE0zhJOlb4M/9ENizGFxl9HF+he/y1yVoYJid+kcesIm7tbHha5yyo40BH8mJxRG
QgGacmfWyW9DSADl39wI5NF4On30V/42x4wX950ALMS7j45FiIJWi7RBTrYgocnM
v3y/N9qNj/86ZE8/ePvAKibgZ+kR9fEUgjhz5dxas4Osgc5x0kE+PEhVH2JybOTm
kWcCD04je54ZyHHsGtj2iNBVeICV/ZsCmlKKEqeHTjC9j9NHH10WqhoeTodzVi+M
v1uamhcARVdqT7/zDwI0xNQW7mx+6A8R8TddGpbo0US4uC+gcYLO6AZHaHWuAHvV
V61pDJ1kWweGZ7UZY66Hh7Z/6wY9Soo8AnYRprrGYlV/KCi/vnOxHYvS0Jp8xpI8
S6Bc5i06pX67T/vdMte9j0o8KhZiIsKDscHJPgQl/tVtt+GJQJO3DyUURhBsLELM
nNHoXmUlqRcklh9CbtGKh5Xb31JYiV5g2579Qn0yAadiuleFalXFO9Bowc7WO79E
dmbmt6oPaZKu342J6IFgSNz99arX5oPpVKGyKKzUAC3An+OoyeFX1UwycRBYqm/p
6oGN7J+K2YdnT1v0awmeQSDR9DcPpCXNMQ9CdbSAm0o4s6d7Kv7d0uwXervMcpKk
WS9AkyyAJqUxu18M/Xp4aNQSTT87Th1i5UZg2ROju4Z9HNYa1quosqcWAXYP40X4
xVNQxhXT7/PLCAIgO4g4Byf5U4wRT5mgcQGOJd4xE7reIBC+TXV+m2qGaO9hOe6e
lYKuejr3qdlr/aqOQyaCB7H+JtXXer/XAhvhbSO4q4SKlWe2WnvrHj+QutMs3YgI
Ib+mksCaDYjFc2q79PenjY1RMNqkUI+UJM8c+DJoak7K42yZteNxSfsbegq/bgbt
b74wRnYTlxOimZO6S37fKSUv9IWmPVPGySf6DX34pdW40AEKvWpF9ZpEjcKoekxk
uwQ5YJIbx3j1C+RmkWcQzxZtc6IRlcaf/Ff8YJ6wqbiROiFAlw5OImQugTn2bnGm
hhN5QzWPE4QbHN5ufKCtwAyFTzdQhMjQl/PexOXo0IoNm5B2tbjxlyYmBKRk5iVu
5gAWJAoNZ/6ODDpmSbbr/ZEzLCFvAZsgwRxZbmC+Fh0OorfMssOvLm83DIvZw530
/MpSeaS9gxbqj16ajmwSnwqTDGjgx0KFAIzEi0z2QWxHfd0dS1tO5BQ0L6gMZSvH
Mt31iy5ev/lsc1dt50NcS61lByLLlKdKYbsupNhUk0zxtHc7Uk0WtOu3/WQjb581
BCrPgi/W7+2G9LxP8r3pUG6ark0NrP18i/zA4AEJLju88iea5P9GHSej8U3Soqsn
uckdZGPMsGURai4cJl8+oDchlHzpWhISA4Cqa4LkdWhpYa6DEn68DTRm4MoPqKRC
FA5sk7Qns3UoCHDym8TFFoMUdx4FRjKkPXdiNp59HknOq8JHJ0xLXBl/xb/Mzems
FPjvMbteIYRB/w4hDrHOejcLNIUhkvNVdTonql1qr+V7RANQihBuhIJrQ3p36gW9
s68zgLwVm5K7hKnCu55vLOWU/qH7bh+fnhOquBLhMZBQw/BW8T7Lv75v9ucQE3QK
XMZe68RBcoZh18PYffgVP49ZvmvulymlRExphM7SBBaporg0nBR8pQD4RxMnIPOJ
GrVS+ux0B6gWptSlfycKJkUNE+uElVagQU2KQ2Vv1Yh4yMuKHulVU89/TXmGXFPD
bJn/pUVLIRMru3FCU+72fAE8zHEOqrDZ3kYl0e7qI/nu0dzATY5Tq2vxRGFg3uLa
+1RVeWoT+gSlY8aqzmnxX0Iipwhvr00TV30bldI2of8aj15nQoIDcOQOmhhNA825
6r7p2uA45/a3LPuhyJRKu94WS22XFit1whR/VXzKlv6X4phOZ3vviX8Bqpv82vgh
QaFgtmnCslPDa5YbduVtRNHOlBk+Syfkp4ux47awTVqBf0KihVB2gCNjMRp0DGkO
0JnHzSadUlyzUm0KypiqGcrK24kL3bdQUwsMdujq5FsEYSbuRw+Bq00FmrD2a1ah
05ztqciDfh/BQd7vg1+HXMyinYnNfEu5gZQ7PUEsPxYJdKOVwyndFOAMSoEZOfOD
uA2H3VDYwcM23W9NO5TKIrvT74sLyoSf3eGRxFJugwX9jvAo4SjWv3Ibyhclt6GH
aytvV6IPWTbUFGI7cSn1br99fYkPym+TQLew+6oVdFi70TquqEmlAPV+DxTf2hJj
nf2DNgYLzPLAjSF6Z3iynyhH5/ib6ZetnM+QdzSNU35vppOOHUwtyFwBf35/U+tk
mQOhzQKy2gEhqoBKVKywIC+c3H6sI4ZCbW5MK9ZyngmtRZ4XQHgAodWLgUWeS0HN
96fayTw1FeuXCxgGOkwFKUcS62WpMetWWTBRhP3cw0u8NvnG9mgiTv5xWQ8YDjzq
WN+D/R2HTCQPFupOF0hM54u3XQef/XSnabmNbORq1/v/Blkbj2wK8okHZWmKeiPx
XWOJVsaRXv1IgXHk4bYhGmZcfQ8HV37TaoHbyMrYVwc/U7243OCNg6vUvh7KegDg
skVhhM6Wwqp/Bv/4K2WGmx8R/93KZuOrvR7J5OqND+QymECWG8mHk2X0rU51rROZ
3C5LIEem2dlm79/WATHmg4RZkU4v0Xw5W+LjW80tOJVhlI/NZzwb6Gp5cyJpVu2z
T583cVH7VsyyUcK3EtcFglG9N2rQkne28IGQEJpnuNTtWtTwbFBuC6hWxM40bWyc
AUhUEsvZmaMKj2DY/GcpSVVqjIDuBiQS2Duptdpyu8FSTbT1Q8hrT7pLvCimChx7
YrE0ORDzm5A3HzUiYGyCHgiIhRQOHdapumf3dJhH9O4rOHtlvyyOKI/iyIJYRElS
CCD7aa+cmAp+yWSFQhnqHPKkEvWtagB1KKNhVnjOquWHjDAGB/DWJ7lPcmqVPF5N
EfbVjbAcdBji6UWca88EV4VYZcA78q46s+h4oHWudvGIF4YT8Lxd2wFwkksY/qF+
08ds0G1PDuV7GjjWMGMBv1vxOSVPRS2sBFkkmPFbnNTDi8kJC5N8EKrIv2MBfm0r
ZRRcr6+DUz5DVBG/So9FzSxpXpwueDQFnr2ZGyOg9V5P85eZV1/6yDy45FZto16t
T4qUfthvPVGlnzl6iEtH40swkozNf9L+9KbB+7OfFWdw/tycqeyGcOlg9wFacPj+
s70vA/phQMc4AyynF8iHtOTJozJB028J6Nnu4kPWAuKHR1UmVWaSaDhObnUN8CO+
gFIKTAyec+/aIGm9Kxxvedv49tkpe+qOWoZwDn7LS9zc3hoZwNkOnSRy9GHKOynP
UyuEhiw9rOd8+R3t6ojgKaH+mL3yVXkww0SNr65NOplzseycG1kGatbqvTiXy9tq
OFOTegtHPGRJ5z97tYijAFrMKfkeWXJZBg54jlAnJz/bntCHFuhqXofPR7XMvFWL
8BJGTZkrdDhNWB6PSpXx+tnS1KJRYFAG/1SEPwaDUVm/n/kEJyRSGS7bAXqIM0Vy
BZYegqgsNnvErscKQRqHu1SpqzZA5CSrdV8p5kUvPUa/QQSzqpjPzst/I1Z6vZHn
KyRUUljoCCC9627ThicAS766RU+WrRkWl/uzN8iZfrCZfiRk7PGK2XLlA+VGnrbj
ykVhrgXxS2mSV2lwz+1JG/rbRk21oxtGhRDTOgpNIxdGuVZI3pekm46vwDLWM5B9
EbtkszACrGMtTxkZ9N8MWF4tMAG12wQKGzX8cc4Q7vYLHkVFqCjfzfnD6ZVMlgzb
0k0/PKAJp15NE4ClJzromaYRSiuwnL135Jyuf/W5A+QKD+bqEzdQ9JMZZtwN/mPb
wI76xQS2RZbvkrki73WRrO/B4UNLqMzjx1wohO7byTir6uOwApGUGlRcFTefkITz
Qpfs88g/AfJlEThIB0nIE96NQEVNTroF3ipKZiHsVaKoLJo14lznAmF8SoLiN53c
TwI6dghYiW9O8HMb4cFGCNTfQaX8ZYzUJA332dn4q0PakMNxt++LIfN6wOWlRJeU
29q3555vEJB0CfuWgffditU4rLkvWn7XIRCvWBdtvGmQQ6PLhgTYB+HBpHUKpX+U
4GCpzFkJcvKYqjc28SzilSJJb80eAzzatlrIra1vf7qqRbHI0pX8B6VG74SoVoKh
psF7qmHE38hr8Vp9BLhsIHs7zV0KnfJKjwMtoTK0VkUY9+30krojwcGw8S6y5zWA
8veRlGjp9atPPwUr59+D22HAFUrwIhhSTsw9dNkqiceAwQqC32BN4HMxIKP7lr85
BNqN+6fTZ90RBtygBcm4WVlrEclY3UG5G4Dx0jLKKqLHJOjmqrd2dpMxJz2usPy9
SDSoEyfUTD/GRvowaccpctfXyNHS8xG/bh8wq4OM3a4pmcyIGnS8imp474nEIPRM
rkzf7oQd15QM3jqGOD48Lr3+npgtTSdDK7p2yRR71bij+aIAxZg3NryK0p3RlF8C
Xh3ADtSn1EZnof9CKqNfTLkmJhcSPunMkGIBh1o929NARxDcWYWyKCkQjuC/DNqG
XFwY2BT//9uuCrAQ9SNGefBcNjjX5YEqR6VLWXxviYvSk8PdON69/jFpV0k7X6GA
XqtFO/2SC8SmHBNFOAeTx8F9CDOoxJK353wFmGLwr8irkw0k1k/9yz7bT69y17R5
IYN2trigipJkBcpEyZGO5HLwjMX8is9xmbBmqRJsPvuPQL4N8MJPx+2PFc+uqUBf
AJd2I8+8wATvaUkizC5d2oyHP3l7PyFeHywhafKWgIaY2jRTEmcfusMySIq0kZ38
deSf70L1kRAKpvqiuFou7J7oyyqHZ+uPuMOA+FHUWtryEBSc3zD+DEpzQ3NC7CCc
7/OL5tsBdE6Mzdok6xmwLa7KEIAr/07udRPlP48I7FaOrNubvq6BuO7FGzJCfOnJ
NyapugkdYk3D0VSq/d8zSisdjDd14ocKriVv6Xr7CVk8VLW7R7k/xHX2xaf7uym7
aNXuAl/vL7nEmc5AQvGTgeM6S6VeC69K6YNcds66NQqJlx2SG+plWD/vFQ/vlSqH
8kkF8SgM9wL5Gc6x32eYiYzD3+64+kksmSSTrGsEqmgNCciO0pnXzUmoNhQ8ruTK
CmGJZpAL5lqqjDsdPPAvrCdtOQxyJxCM5S/TQRjRySunvCtlFFtbQL/TyNvwSFCy
Fsr/bfUop1CDc4akIctpGQFyVGpu/jrLXCv7L7j5xsO+PDfy9qjWvuLje3zgUCtI
+WbPqP9Xt5dbPGmxkYFtRqKXXPfekzHLuYTN+mRgET7Wga8owKJn0WUpWkHqmVEl
Ev8nN64xK4DBfLjSJH/4xLqok1UFJ/Xr/K3gA9d0PNmaB02e2qnUttEgXBQqUGhR
J5ehU7zXMKaQqZYA5OhBO3W74sLcdfybGhNfGokGJqrKjx+oKQ2BjVnRzB54AX1J
07irQddosvC6LTPZv1UlqgToEnkpVxJBETPw3xtZN+S8SRtUEJMJpO7PSTi/9IR9
a20cy4bb/wq5NXKs0hwkkFwc4jYc9dGSl78hSrvHt00oaQRR71fo5tMG3caiVVxz
qmjEcYZ+14Jfv97a+6NXNKuvAN3lf8odO20jdM9UN8KSVAoqhM8fQuu0xMA9Ekas
f38aWw5QI1XI5DZl6DGnKFVkSOnon6S0GILsSOz+Z3omiB3tZDhdgmqupkrSNKFN
d8jpxIj0qf5lD8j2n78QCOgFpTLr5aoA8Vuu+KLQpfWm1rFiFIhy7ENfymRDgwGV
0iG05VSObS0Mpc2ASvxKfusaJptLMs/b+mgoEJZx7jjbmYHkkiiXY36dZEX1OB5E
o7l5UA1NPuPKII99k9AoAkPPjvpM1q6kbJoVWaSyX3aqbMXgAZ+dFEYWRgfWkXzp
Ns4HpVsVtrvDWyVzgCpiq8rHZ3qS0tzr7iWSbidEdB1rhPHfN12oqRB5W9lw6xoY
SkQjO7iMyMS7rPSclrGvp55Q0lhJRXcDSJRsVlPosXe0H0vWpXdCiqIJUJcOmZzC
2xR6u8WJuaon8ITE1V9pgYqGssqqwmzISCmci6djByqrtDyG/4urwQ3mTwNwR5jT
V3rzcfn4/nzs/myA/UkDhbxIv8o+T+y2lgIz51Kj0xwuV2SYhUxkXwR33GrECbWg
mSUUQ9dAaadFWMxOCB70ogKOyVcY4vL7YZ1ZV8y3UOCjQFetvpFExe3pAMlM6gHa
rCbvMIOfsgcEiYgtBdA5X5taBpJwH1rQgvPGDvv7q+dws8/nbMdRdquB2Qx8FRxA
sPp1oCihhuqxj2knpUgCdtUMrWQOe1MC6HyC7fM/slpfSOpb/RR6ZRBHBH/fnSOw
FxRzHIdwaC1K9Ztprt7noDzA4xpT0o07f6aTnsO+G5K6GfQIXklau0C2OLIRov4K
Wm1b735uctjFWuuWQxTr5X0vxSuxsbmyHhQ05twctqlHbZkVt45ElpwIilu29j8h
pnbGuJfdGOfOKxIz4WHccqfydR4AQqS+Qf62IwwQ0FG3Xv9HnmZcln+G6zdIzaiy
atAnaOaMI+5LmKQbmXKOfhidFEF9VLYbinHTF0VtPsdo0xZYhBhSL/kFdaQLwubh
g0vUpBEAtBhG/8y43LBUYTpKdJWBqYJxxaKidPb6pobpMOrlkZzj1oVrpJEPKLoW
3rFSp/ZvQQbT+9hMC03ae11Jw++YRxi1ywyAJJzbdWjpR8Y4rgVyIV9q4jMoQRpv
zZohCeYOMVcPMcQAelTqeF7CGV9vem0ACVjbnsKLRaaWR4ig/gj30U1ml0lu8zKA
KSeKrlO0SCd0KbK8sZe1Omp055xLoVt7wEK1UuX/nvzIJSvz4O0sj+hTm29HKcQl
zVNy9Es8M/zjlcoTFjDicVBpIEv1Hmw+kAvSDl0djYCDBGC+mP6+xHjyXK9Tvm1k
4d3r6ajQoiQRIH/x6UV9MLsscz92KSaxMXaD0f+PK+hv95q3S1fyP7DEbHf6CLEO
8ienqc++rwX0riSEYmadf6sUwccVkDHOPuIXOd1GGmehHfus7njsdsqzA/kqLd7M
YVQlbU6+QeaNbsZeE1M6WwMi5/6M6SPonPcpy6KDslP3V1L2nX/6il4AXV/rLhwh
pYgswq9fqYs/AXcYShHeEpRZKb8UFCUQH8witbTRDCc2BRp8riTrfUD0Kp2w6dhI
DlT4wH9HWp/5TXTw5gTuNVAxb1TJFxrmJcCrxwfuanSDgQ9SgxaLtgeTEfaeR9x1
qe/2wPKCXODQE1RN9Vf61yeZgYHQ6yODJA5Tyato46Nh+eP+OUMcqh+h6rOqqSVK
9mvlSPrUd1GlrFS3bOFjJSLPoc2PYUSxKT/hlZ7WQB2kuctpcaWb/uI6DYHE16St
cvuUUutWjNODV6qyOYCOSCZva7rgySKjI4x5LpT6hB75rF/BarN5eht4o6FT7YLc
0OCoV/C4CmRSorPIvCHuR3uPF3N9QZODwdt8puKolIQwVjuDJ78M3ZTjo8EBAVB6
5OEz+9ImZFjJtAVjOuwGs/me87LdctIbQUNbbglKXqzbg0yEUsdGoQbpNpIO2MXr
SNKi8lj3otepvAKqHDv05a1e2Z4U2qZngRnX8NASZ1lNvYC7mZg7jgCKzxARmUX4
plORPZQvPTx0/v86ESXwy/jLFtFnV5qc4MHXdRJwNm8a75ToSP9vrC/fz4Kc+jya
/o7m7TEzf7kMib0ZRURT6pFXzgyFXej5RzXa47/lOx2jDGqVn6ZgHRyv8W5sisrw
9SpKSLlM9VewVqnMLkW45ishUJxl69ZllttqGlEWuGnfsAXFbkbZmIfLM25pmZSI
9hhPXDwGM9gGoPNB5ra8LkiKAv5gB5kTMr835PksGvmtJqtSP/s907ng5gBNlB6D
mVCwtODFS8Z/foFL+WqVMjiWkbOHNMzrSnVWqPARWpNeqxoQPzu1FwW2o6KMirfK
JvBlWHyiyVDZUOqfCCYDvP07FxC/uBKBsXKXMzDtFQb70hUA9tp1H7+x3GIR5llM
3nzdS7JjbHmyZ5VT3Fo4T2oE2Qvu5eE/jtdU7TJxoyo/98HqJUIgNbNw3Odf0/n5
4IdGkwLZieemiAYJvtkT3Xw5cG6OLG9n5UCQ+Qsbi80AyNN/UpFymvAnnJJo8ZjK
t9K8xfh8kyIfQ8z799oCtCaVrMpMf/fXu381LWa9iOt43gWR3XxVB0OMr3Mmr4sG
lWni5phgmu6zx2PrHPXrDGEtYJADqxQicpE1pnFNIOGze5+XMGTgRm544+M847fu
PLMR7hsUC6ELEMoVq3ICe8yhQe4BCusExeTvniUtDlvdXnxw43fYDpUpW0iQpXU0
rUxX0yK0ke8ZoVK45C3vtKhYxeYl+YAITqTYA2s3cx1BChbPxkug7o/ruUqPQKwS
Jpf9iIPPQdrKQ/BPmHMMcqJ1NpNG9MYbt2LtSx60HhIOJxuxs6xoqo58i71+OHQ5
+5Eld2PKekes64BBY5Rbpe70B2wSDAKSHaZ/9KqvnxrtxjUydNnkb9kM3IhtDld+
KIhBgnAilbaEPlpSq3Z1S1lQgSRoLF+dzP633pUKCRttRQYJqkws7N6dL4UuQQAr
u71ytwBrKeL0nU2/dJPyM7ykXQ1AvUCQA09STAOBSTw1YJ0xFasQd2Ugwkh/8/t+
D/fg8z4iwdnxwooTE1awK1ie98tYZmGXXlq+E19b1BtT/ioHLiDA/qRdMZeTwmpz
FugKwP/b7iXOL8XTd2qWpOEuNWYunrTfYijE7X3t18NJWAaeh33lX2AFqe5ajg3w
dZ+wmvhHABmI7SgjPAZH9UcYhN3GeuaD0noxUM4OfYrdzlU3hCSHCPre8+AF+c/J
59jBhjqQZgS1uclzkeOeRFcPcI2Vcpms1zsumdWXcAJop+If1km3gTOJdGpd75Fa
HwD3m6wMVhLUSiqTuLq75civrEtgJKY0hGVGtuKWJ+xKCUmtkM4S/W24PzjM0+Gq
bKW89f5d2uyFwQ2jWUGiLHFt1PgCT9bsi9Lr7wBmSSxaXZnQ2wqKuwB251rN28L8
kH7GIuzCAeDJNCo831IP2/EWkRWkeIS2o4zy/igbLoewfg1hp5qhmg7gAF4jUUfE
jhqYdk1CL3xdvt/V3e0ldV/VX05mUoraiOtbZMj/ZHd89RJlJ3BlTI8I9SUHxjnM
LfG015lpYJAq2YEeB9S3hiwZ3M7LVy03/Wq1P8Z1KXiNKlRDHxi7+5sFuXmaSZLO
KGfXqnFk7J37rm+ia5LGg1kObRpTJS+xerKWmklmp8xEP9IA2vIxzcXoUz25OCmU
YM2r2r2uphECjxusrsWUEt8f7kwq+JDf7rD85lfLUgJBfLw/bnFjlVIywVhaAk8A
l/5p9WEeL4VEHh11OBQywtbEzZA8PhHmIzpJ62oWRVO0iWAvJiknrude+Aqqy0F0
rhYFRA9gelk7rlxHA1WrQcTwoCkHXpgybOoGW44MvVHyUVCOWZz4ijqQkj4QN2z5
0FWT4LF1shPcmxEfHI6UyagoORouu4/69ixl79G/WKIp+JCE/J7J+NSEVxU+Daa2
vQrm7Gw6/QYA1uHTEDKzeOr2km9ADSq59DCLfRwaf7zdJCwhraS8CZiFNTfzuWtT
uG6oKqGaZHGdNA59kmlY1zgHimAUkd4WKCdxGfLVJJz9/GyVczbSPOEXUO5XmQhT
WIrvHCYyZUNA69e0Tu8VeBcwnZbvOd6c4vVgRsoLf8bVlHgaA+Ld2nzXAJntixpM
F4S7ZUlLfltlBxOMXraK/v3++VOUROVSJCfjTpzvNAlMmaRzeHmruCmK6OC5/l+B
RdzdeRwr+Z1Netl4OO+yNQ3XN2zEOlvDLgV2IcMoQ9cjHpuEAoo5Nn8/93X8uwbR
qaX2oVHPFmX5hH92pHU//gafWz8fYVrgf7O+BzaNC57cC+Vi1J5gIE94e6gXK4my
aGWKzLFfpkQ8jSCz6ljcUoePnqY8QYBd4vjAoU+Q0dsGLpNP2TbxcGpuTJRKl5Zq
MilU20Em1++ZlzgFnVUDWlOzXTIu1V7bPscl00ZoGuxmwwd5ypHeV8eqpxfW5ddl
PHfXC+lhJblp+sDSJYxDJrGK63qyPA4PFPTK31aERkJ0wWlfwAWxbFTaKamqR+i0
cQg9XOZ5yStjQTRJIMY1CTUxWR26+2FMkuxlZXHBk3CeL8LoGFcPf1DA/N6ZQZYU
UjvJprdxkonouIV99zp2A3PltwoDK0jBYD3smLh/lvQhv7qx4Rs/c0qSo4dKifaw
tPKtxLuDTQ0G15VC44G+BnuY4+BkqDFa4yFKRl2UCrY2APcJF3FdgJloDst3o8qZ
gNb9eIBdjxDs9QwAzevw1Y36LebrwD0Pv/sEdlhuIOwWw+R+9z3ScX8rH363JJFV
sY9/743YXzW8Tgu2hlZh4CXkYdc8p4zoIp989nJTYuSP6mjJfxkILfkfp6FyHeHl
j3xRwUxWlz0kuI06KY7NCurNOXAf5Vn2rysoszrIUKQhwN8yr6EOYSalAqz4fiTm
oFSTCiPhyPDi7opwgfLzJikzrUN8i3XYjry8vjCE9+x6gTp3gaupFCAXywa47ew+
+4979+vJjNbEAgfnqvZkXwIxPrfcm2YH0G7xvm5V7UGSQDjaV7ee5y0qTRzXKWx5
Bp/EwXwWuD6agUv6ZoigLZsKyJjAQMGnCvPG1VfPCeyP2JU77W3Qo9Q0qg5k9ill
UjBe1dXOO5DgFfmUzDntz89Y3jK12XsZzXi5TmiYdUrnMHUVxbqOOlpPEA2VkNMH
k2MtN/gRUfJFWdtBMZ2uiljTjguDbogu/uPqBHPJ80Rnf6O1bk5pzu+nLiq0J8BX
mJSA8/fDutMGnQ+8Rn/0WK1Q3cItR2P4UMLXWpGBZtM1Qvuo/fAnOBB+GsQsv5Hi
irh6tN9wapCK+8dz4VqhR94RIcUnHVTj4R+8mlp+tys8MS/VI4nbU9OfARjVXkJU
mwY9QXoww8GH1bCD+wPIJf6+R/tYex9WhSWwoH3x74Cwz7PHuxe84B9Jxe3PpZff
0opYSa9cAHqYqQvGsg3jpSQg8WINRBVOElwJHaaqSeEoBXs+qeuBJmAUZEmDLO7A
Ezs71iBMdxYvE2dc5BFXo/kZNMCtXJ2T4aqm2wy2u7D+ZZCRCptjfXp9k27ibgq2
NvNoxZuPmRk98suH/+KlUsrNWdNa00exIGmLbhbSaCu8NNyLS2g36Rx3NR9EKmwK
Zxom+Gp9wufQk9rblzn/k08/fw0tof4/bRMDTS9Ush68bJAj0twN4nCPDP9pui6e
1Sz90tAvOW1Gietg4Go86xd3O6+Li2p7R2Q90Rw07Dn/OiFog/WF7ia+AYUSuULK
gVBY1sjZldq9uCOzSzBz6/p++mq+1YhjHau61lLJtvRfevT8/IeE8wZdnIeF3r3Z
V82saLEAUu4LLBjbZyHLyEpaPkF0R8/FoEBozR8gqvqaEKZm0g1yLH33rZljexD1
IxYaA1tYnybB5OzOmltX/lEDKaDZtbwEj8ZG4kav8djwJQqZwQz3XuZYiSvjYCMs
lpW+HYfz6Rg9Q2/C3JjUr3JQjkOFfxEt2ue3ZwkrG2Bmz0HhmTIGO5rKLWRRk4xH
B8WBHuqaKz9xeIpOMoOIA2LV7ZpB1LaGI8xLs+Kgix4R/uxWJz7XQqphB9ZpmqMx
LgAdgnqxCdctkw+ITxhWe2pkl3S1ZRJHCFO+bPHsqySwtws1WS8IICa/cQf2DdiE
PkxdInLZ3OIvDrV0ORBobuz2tXZAPB+tvqD4XeIpFzzbQVzUVcjdjg0XK9f2qr3u
QhXyZdA0za9VmBeH92wBg7m/wOMQ8/YkB3a1HUqQQZNgMbofXRixS/IwhqZhdJgJ
CZwX1/ck1zU4ItDPacmMW94lrYdBlbucS7SCUcQx3KDAWF6EyvMxNQpu8egUKdUV
+bd+J/e4xCip5m6/gxhQA9bfcaGJI1OaYovyCIxavpu7ohbfmv8+WRHcNIcN2NO9
QhOT+zZfOhNNQs34qQelVGAOTzRxiSjjyAygOsrXRqrpxlY7nG8MYlqUTaLDFsbZ
lmMszTQ33qRrXJ7zIatpwtLSGUkQIvFoognTFUf64X8rZhhROUjt1hKZYDdzBCRj
hALHVhRIGuvmkTSgTemyyR2Awn8rGxioqkdi+0RuPWsF6r01qtg8UlrliHrLKjX9
RAxrGF8wZEWHkjRIrJBF41nQh+/R3XPW7nRqUTbMOVnoAi+4ksQWdus4vGO6vBKl
hppPKOT7wgUYuulcF62G9fEHBVZG5ReQHRYlVxmkI5xdPK39HQWZhh6lfUDv6zjA
5Elzxnl5bprgLZ1EXmAJpKlqHl8acGc6rckH5gzAOpW66yvbhvvmTNVtcHIMeyYa
GFZltr9uTekUgIpHERrYYiN5Z5jPddJAcOenpO5bduf6RsQeE+UJZNePi67R+VKD
yIOCKcCDNMltO+plq2LAomDximHxiUYJP7rxqcP+wGNtcJAWysmgI1KPcC8sn306
uZts7brZo08t1TGs7Bkw+mEnjVOaVmLSqtfHs03+a91ExdcJlmp7SWdY7rrl4Z/L
eGN8IoRmNNKS0ZIyyE9ruZroReezSTdcjSmU2i+rSXayzf/+v/we3ma9iuu7XTEc
WhCkkyBJEEj/33TmBM6u41SpffVWoUWErfsCmrqGRRSv475MkSqHRss4Rdd//kPy
N9LYkTSIN3tS8eiiQMhkn4RwWiJypaMpUshdVteBQq78jXgKXLxQ6U76xmyvVbqx
ntl1jOrilRivtazCN5nBqtgyUELAHlpOSmhaDkQf/49Ml2glOxP6y5QocNOAkT7Z
NjKkPoYLev7q1grFJ5TVam/2Ks6dJXOWgb7aeDYEYSCo5UxFHDjo2wCesT61Y4sJ
gKQvJdVakQmn62WqzRU7Rcpxw9on2CfAw0gJ/+rjF2cd4hILFcCHfmyaplIjI4QL
5UEmeX0NTRUBHGhZrmGcb9VPkzv/xaDg3vkMDjTs3bE9im0DpK2wMYesbQgp+I7v
rZaDCuN/xxTypQdh7rwfAkaJcGfULE7Doxy4hNZntai2oMjmktdLp6XKG2I+uYb0
DgwOBP/o4O8jbZHmDKziNufBuXi46fNJVLqJSnuSdR2esNDifWk5EHHxZJJg+gkT
8tvumkX22w7IUKqZ2FOkRegMu47BSMUY3PTuU0fU9SHmEWYWiboOZDSDTM54FDe9
aNht1x2Q3rDb8/YhJLlYd7a//WxAq1NnOXo4ppsa3xDdVBRLajWRWZmuf+Z5Yg+C
bAPwJu3qAiU6abhOg7CCFAOq5+TYfRxloAjQcI167e3fOleUKdLYq0RyjQ8g8hjM
r3MPpHlgscXnil6sazuW493zXa2utAQ/LsY9AylEEAH4rU5CB0HQY1knLS45Vo5L
t+zbGdaoQ5Enxb5A6ACrDWenwkILwys2Uax37Psp7g/V7ZVSSCa0Kf2Gd9OJWOW8
yvulQnbsjbZ6IBbpvUzZvNlbSwXx1PwHXQ/86vH3wYrLmOLRbiSBuBUsgk+tawuB
j3zO7WnRipd4IW4mXNOoIeu4K4EovomCCnFk83+OZbduMOwQlT1PjnJFU5rs2RpF
HhyDnx9NgdlJ1eFxcUFS0OmlqtjC5c4s95NhrYs5itV84RtR8CQZbv49o7BNyVB7
kxN+eGeV0e1pOmRD9hdSop++3/uljh55tgJRuIprtq09+ybiiBBXgeSujBZ4NU1a
FL0AJ3Dqb3oy2X7BW8TSoE73TOtINxoUlYOE2PRlBa7OABqXzpzWZUaLfs966TgZ
jduSzpqvJZ8xTdZ4wwYhm6UnOV12LCUqTwfOr1wuBupVIbfwyQwzY/DErJfKh6Oy
Drwb1vie8XwLeME7My+a8VlZtJLcafD9xhokd2ghUksch0ZNtqaEPu1vIzlWikRs
DsegxGWaICK8hjMLi2KV6sB3Of8PH7wIFy1TBLU6aPckqW659Rmy4gQJlXXqvie7
8cclcJVTXu8p5LW1L681MYpo13hTTJvu/jVUYTbV6AmdyZWleFHOQdVDAIN5PEK2
jZ8wLmy/x93EXEkFXjYYVyFjkaDZwwTKksxPw+n/l/AH3Fq2KlAXEb/gpn2FCh2n
t67isQ/39dqHRq6CbyNyyclPq5ymIA8ETK2YAKzB88ESGpmICKEWnIlXV3tx+EKf
+aMUDSNGqUDM95PkSnUZsKCjwNw+zudMziAmfZ8G9ns0Pb/0OdZTMzBzhUZBW5C2
A5ZpWGQLhrCA9skhJ4lLRxzRWD5KLqSKwFeJsvP+5e02IJA4uaRGf43HIGl39URb
nfDaF3e6+H5sRyalP6FlYTIY7ofa5iC5c5HO7GRzTy1neUeralbl5avD5bTB1Hqc
7Mr9ZvSUb0WWlfanUXI19WNstzCvZEsFguUn2XxUA7QqCU6ZCOj8cFWsIR90Bmy8
G7RzOWGp7Ho8gtQeTY4eu+rZm0ZafBgGPjiS4plFqHakfam+LVe3G0mkgInQsj8i
9jRVcunZVQ2PyfCGKD52TSyN3pX/3Rtm0C9NebQxGh2I+LaOnfkQuhQrH3io22BV
jDC72dg3syyKNp/Xa1P2p8y4pHOZWPcJCyMMM2YeilnJ5Rn8EbBFoH5syln3TN1Z
lh9LOB6dTFIzl6uP3eo9thiX9KnaBjkD6Mu6YUxmTXR328yGb6CrY1ZYlUonn7yg
A9ZTgsfCinFVefNovgZlNtN1aeqvFfeCxrKkFX2ixyq2Yf32yLKcOdm03vMf9aiQ
4GkixZ8PM/WMXLQGBaV7hLgyHPbQsz/vBDjPvzvpnezWROS8xibRxG2wOjknN0qB
GZBGUQ7jAn/heMYUkej096Oio0SwM1Ees6XhK15DTBUq8FAvUbujUEXO71ii/MiQ
PFs0pS1e7gGZU7GoZby//HIcKQ6faMCi9sZRma9fvQ3rIF30mlCj/NtdnSswqlrt
jult9VFQRZ1P/JTw5gsL2DT8CvEBprg7oIe5WlEM0KtraTJGlqL+7+aZWOg206xT
HiDYo1O04z0T1Nfygj2LMvzyLIZCrDc5ZjVUbXt76NUNiOH4vhm/Ay3Kp4t8HCQN
Md7w28hpwH+7xRRULS0Vk9XniN+81tM7QWgS7IzeYhN0Os4uWLIJaG8yrq7GiH7E
hb5Q05p8qo3qwO0N3NRZTKgS478FSvTstMgX6GYvumPanQmnsBytDXaTHLi+RZZw
b+vL98OmNlBi+lq4R/HTVPj3S9uTe6AB8Uws+XtXriawx4XMNgNZo5a2xLndRGn0
5fx+RqBZs4CKfF6H0EQ3Eu+exMry3MyF2C5uCrmJ5MK4NIlvyZ+Aq93YtcecZ0WH
A2mjX1RV74bwQfRXm+Frx0i25hmNCRDTqHw6OFnP8kKNEAvgIMKaBis9R4SFrhaN
lycC/u4cO77oOOhGbnfiQyWAgZvXcetaP/HDiYN1+QkUPDee3pzIArSiEC50rYIE
hJZdqRiiiqEcodeKmwQvV8r95LDJWYnuq2N/aj1A0CmSMtQrN7V6Bdv4IrNXUXQ0
+QehFZ39SR0HedvTB2J2Jyh4/ulKIDV1CCDLQ4UDQ0bjOCliKSP3UPB+Sp+AAL7y
S/irN1gG3dE1c0JqVMvY7QlyzTzXV65E6bQHNnpbMi5PvipV6pqLTkoKv4bnI3XZ
1146v6nlk3syhwHWX6BJeChl91hi/psXEh8DDyhqX2m79MAFHHrxtDuW2RzeBwvI
ISYtZ3rxwV9Bpc8xgfNwr+lij87UKMS3ESdzk3+T4u0w8ffP1iYe7ZNlEjuthfSI
tmr0PIKbwUoJH3Hh3bS76btt2pvGuyI5Kj+pO3GFw6ZASv5i+GVdbhqEHVi66DO6
5rObm6KMiW+2pj4Z6Fo5rZW10MhmyQl5x5cioFsZij+mrPHkLLlHzIW8zJx33cv9
bne+j3oDl/VNcvUKfz+HAZVtr6406XTEP5/Iretl7Al/4ubcS6z6F1vVnh2nD4wg
HWEg/nZ3+/eEsj2MBN1p6hQdalqijLJFI6Kr5fY71uMJqYH3OxaNK0Kz1lgP+fh4
TjKmsn6DYJu87rlK9UoWap/tRNOvVLIFYxCu8IE4aP9i9Lv1UCdhaxta4GSjYWao
/galsst8QBfHoUl3r8i1tLIuFfN2ww8ThgapbL7gbLtokDZT2k473RLlg1LJF4EF
rYJVwuUiW/F+Vrp2FZpf1InCFbhJQPF2SelAZ5wVJ6jBNqQoQ1vHYka/SrUhb+X6
TePW3fk1OAmyR5J1whwDDcy4/ovjk+iAGzEX0G+AM/LYwBEW1XJCu6+GqZjTfp66
bfhIrycjOW/DY+pGUP2vI3lVHhimdpMjVTneH8Grbe11/1wWl3VmKaSUEeZ+DUap
tpLpaxAQ4L+I6lswjTVk+n0F/tMyEoje1krvXhJ8Fcd1Cq3kZhn8r/I6rrPHfiJa
WHMhzOuRfL3u0r98r69oDxKDKkKbwoGsB+L2nBhVaEgPRtXxy4MbdxA7/9et/0M5
dpC+wYeStCcq1EYCQ+dSYjiFwjCerYRUmdAa888LdrP5631gs/nCBrPzXaX4p1n7
mnDennOC+5ZB0WRuNbth5PvAuOsAQTv253lnLd/yZmq+FO3mFVkrWJ0y0ySe2RHo
uoeoDvmNPkEzn73mQPdVLWw81p6wsVYqBeiW0t67Wp53R6vkp2OAYFa6Y5oiv++y
SoDZ1NmwGHk5ApUYg1a5VssEokhj61gkqswZxKzbJsZU+X5bF37HLJyt+dTXjQkD
f+EXIKMan786SUqmN4B4WOfV7Dx0MfL6SpnpS83RfJHJLC3FTVpT9t4iOb/7QPjF
NRaXvfuAy1SKjQW5P+FPEtfX7Fr5NsWeAwiGrL5Z0HoM4sMf4tJdkpiPwoLRUetN
dALOZCTko0tNFCkZFwj2f7qJ+lJmWY8Ts1F6opgoxq2lDOCLvj7kVh6YHNsKdJA3
ClB/wy/f3wB6soKd/KRl9NQYaRYLMEm8Wp2QRXtw+58l0tTy1ztWJZWHN2rO6Jcc
3FangqGNAsoWXlRcSD/ExXZBKmydxqGLDZiTSvyhunASbJs8PL/Zt/pTvu47N14T
/aaf4PDL6DkgUi4nhu59dprDHJRO33r7B8Jk+SVQOMHy+6998n9TAGQu/jmh21EQ
nsU+F+mlMMsREKlhNBzuuGsJI7t/yiLURjpzlHVEK1dho1iWGsaZ7AHgYr4pdHGQ
/VZF4e4A8f9wMzZbw1g5cXDtWbWJ1aJ8nvsvYO29bR8ghjyMDKIKqrS1ykJydeAt
rF2ZKylr5ettsy+IL/OtaUIZznlHptV4DP6Vw9jIOVDKE/kmEMeUW4gQwTbnVS2G
B6HDUkzbpbuBnPqT0jA7cfFthBh9LhdmUGirDRih7gVn8KFZj/HlYXmqnP7iWlIT
lKXzT/SUtMM7EOBPQ1LUR3bWimTtuovX5q09Io5mguXTJTllGFjCGLg1WbhYU/IR
oEKuXAbDKN9KuEtxZv9k/hJJpHaBrthCR3eDnPTHtKHay1/N3aHEEZcQsYkw8v5d
jjJbX7RYtOHs6xgSmTNmOGGMsJZ6I2SVI9VWRrtWPqXmLyqpvI5BvXd7Qj5N1Uyn
Y+UHNAzT1tyloohl7GlrN74UuN8i6rGUpDaNPL/plts/L4iBU4C4jDxI4gip6c4O
FOJgy6gi/iL5Of5HzFY0Zvysu9i/qgH3myYFH8/Ie5gNd7pf7xc2m8VCGnHxiQad
b4WLPD0m1jyPFLxP+Fku3TRB3pFFxWo7S+oB1ZmmIXcOtcB3uo4u+86Sbb7xC6xw
JnUiZ0K4Oxbk2YQkS6NoOLYb95inDNpsFMhJJ5lfLyXN9R8Gk62LfqZoLcU5mGX2
z+uYoR7PhTPWUI3orWFH/BMiJ5KE2GdTtmT1svLBiNw36uaN5K+S4FraFRjbXYj8
Nb2KOJtgpLKZmguhnrY9U3qz+KomPn1RxDjN8IZ01eBhLyUUq5kkc8K6viC3+Xi8
d2pt8CY3zeUw0166GDZGgUETj5afdbpkgwGj2Sj2RtZS+XjDayd5YXamiPVP/BLE
FbqJXqh+9cg4koxqDoNZVUXiNLjQ5Fws8THyLcsa2HxaaSCT2qNoSCuH/q4Jkirq
9nuA2kQe/BhBaz89K6pqZlXOzbVFGX3o2FbQxbGXevHqqZrPWnpGGhz30MeZwjG3
FGNq//IJ0CP5Pi0RzO6DURT7j4ks7DRHj+gX51ybSXVoZslTaINoY2orrqgJWf6J
C3BICWthLqGjcIzakhszV5AyXDfqttU4LU1GbLzktzPe50rG9XP70ow/NNBL2R4x
StykaWzysV/JBUgTSQDGvkRO+ly0vl//kv7cAZV/o9KfSwdTBz4ecMDDqQolA33d
vTVaoBFSyYIUYSVzTRm+z3z0SIhC8WSy+iYOrlNpwOCrsQ6hrwr3eQHKO4pXzUT9
CTjz/iYu78eUlTn0ZcSaN0S2s17RvrN2/cvoYd4E5iwyxS+MEMxRFpTSoCpHFiFK
/wJ7A7JQwyL4jU2pUueCVlvEHK1Bm9qxFyzaxp/ptxT/z1zIFFXH+h92A2/ekUn7
3BxoacrXLGmujaPg/cXARV4VTnhdmEbJyjjAGNAvOKyVlBMyMPnbWUZSqVCK8rNR
4EohRcyGhvOecJGYgh1AzNl1QGQJ20eHTW0oj4pr+H+QcAUWVt5UoC1xNf9uEYCq
GsxQ7FTZDjQNIfEKW+qMA+f/wHNHyStIYifhR0TsYA5TwRPJUM3BvZ6Zqjo1RpII
GI6SFKGOjFPr/jUsATkScgZ6wyLd3FQO8bPiue/RSaoXaf6gXkY+fZ3s1WW9qp+q
UjqsD+sj6S+el5jr8nXApyZqRiuXOMmn+D1YADRqkf7Yd9huHCT4NEJau9Rrf8+i
1u6tR4U2cZNaUSUru9QbqzlYoUBAuozwAJQ9Y2ovq/lgJo803KgIZ2qXCkpdTAeh
1i1dxnOGAoNDjBDTPKWL3QEztOOLr/Yuf2zWZMiubesfywUd7SPgtSYKLuryNL+P
ndTTB4sQQPN2rb5MTNMvRSpOtxcONQQZBqeF1+0BhfbiW4qXah912FnIGN5o2zdF
Fe7TxugHi6J+x/1ZMvlpUpkKFhzTzm9TjRVwtG6mg7DH1Y1zV+b7SNWxSWeP1Ru0
AnTODkt7oymzuSJC4FeMzhX0l9SyJpq7PxRYPwovjkshxrlOhHKlE2jHf2xpND9z
HzGlYIZ4SaHMXvn3cS87frrJLSQM7FbjBHMWb4ojkxj8+95l9zO3pzMYJpK6y29P
GH/ybHqv3Wp+TgSYh7RukFIbL//rzILvGGKKXJ8Sp+Ea1vNVp+aTgSCRoVpQ9L7Q
0nCr9T1GSdfXtUwdkN92f65ol8dcdu79Ed4dJBazwpzKpUsLVRdW7j7oqxehhJw9
+arhVv+QRkK/HggeLzqrEH47gmXWFp/fP/FmDaY/FJT+Ep5E1Skq5OAiVY4OfmYP
r7VKypYAY5VZLkHlnHpBUQBg576V4TeZk4z/lvvFxnniVOqpTSoCVB8GkXqCj/Mc
Io4nCpkww0KzBfJ8+MbClWYyB5S33lJxrE5hCufY7naiXMFtSPq0hg48bUndWKwR
dOs3jJ+PxtQ0igNc7WeyQVZDP2T8Tr7EzgBzRBOmTBbMTcdQfspYFy4YEuWDfwvX
jfvKlVo6h9GlEKdppbDKvHOgnlG2vS5iv/3/anjoC8Lz7Ab/mfk2uoqW+CtdGwiw
68St5FcJV+g8NK/NAV8fc3pAbsftsKfpWDKoElmhRoHiBOffN3SEE6NHIxfvYKQo
Z0Kkvo4bp6CznMVBC40hjO/uhhCABwfbPrrUTMKljLxzOSRP99l8eB7m1+OAbCLy
l9PNBMFhX0xHUboHU0fTGvlmizfV58ChdsGJj1rQSZCyDsflafTtLnOMdbZa5HSt
j9wCHR7aWD0ARcywekzbw3oXxOj/qlnmgSb7kt+CYQ/vxr33KxRD3NpiT4G9Ea/4
r7MzlSDP2+l4BBKeD4h02T60y7Ca/vO0IouJtknBMAm6NA5xH6dyNzhPIZ4ZwkC+
2Qj8nBW8PEoMp9AtMarpaqy+lpTQZRD05iG9JeBmoVYr6Gig8p4PwpzvLLnJ/+6N
EIXXClG8W7xtIN/MHddXy+PUWMfn8j5V5VtMJo5uI5cl5fo+pGelnOmEozu+Ya6/
DcxOmOu+PvbWYBLLVrcJrtKVM2gHNJOKBdWUduUgXuw0WYSaGVIsWAAFhIgjXGwh
z1+AJBcwnyZgRezR1k/Clm9kuDywBCR/nOThtIqUxnXEzvD2eKaI291GKJtFP8jb
Q2ec8VJWNZnZd70DW6guZQY9fXucXXLOOq5tCc6801FwMzaAwtSES8BWLnshrWWr
oqdmO/lkhEaFqXaTHmFc6UULR+p83c+YelKBr28M8i6tk/lFEecrmb42nc9E/HNH
crRAZUrVAWgu3zmMbDYploRbrahSiaCKoXsMR8HFfL5OPkk48c6DUes3gKDZeEPr
FDqMp2FmWqFN7fEizrHzVoeiE+Ce9/EPuy2dxdLPecJVoWegO3jMqzkCg6FwLeOl
AlIXtlLXyMdM6UOv2m7dcrwBPijQVT0/5pMyOZSdHMzqBwOd25ni+BwePCUqR44u
Slt2Jex8R1t5GSF4yaMBWqn6u3u3W8Z79nJ8ExTmvdDmc9P1dk21nSjY/lP1zDQ2
Icc3Vm6+Q4NI+fjYhl2fSHslFe59+GtzW1cUMry5bDxnaFEmLNwGpeem6xnx1Arj
juj8XR5ha6Cr+c9xmnij7vUO8CPA94hxPkzUG+CGO558XpKchYM2oDHPd8vi5+N/
BOxN4dxdPD5sA7xOkwBbOk315dXHTlpOLZgyq/buHzVTaym++3EH/9JWtvo1RnX2
GZlPXgun0Ce0SrPexDSoPm0poonAQnHtsuf0X0Oy4bD6fokPPEqWRX+01wsduPPz
Wx+qshIw87e/5mSiJq0yOzI6KhaClPidXFgm2nTYpYMijRjrPPaQRYjm84cLA4zU
kGpZuxQw/Iej7ZvK4apIVQWLKq4KNsbWCCoSqI2lrFAPCpc6YdWbqTW/T81fp/uq
CX/9BHo3imud40CT8AIwxI32SpZcUv9K2qFsxb/1+gUfcVB19Og1yJOTOCQaWh9F
Qhzew4IZh5nxhAoRCfsQqUnynFuAxBS3utgvK7c0ZUgrmG1MnT82hHm/gL8p/7Jf
1Cj8skZg3PSK1wbN779DsNysMecPsyJW5iImxnraff+eSzHOqdo+7MpEZigG77Y2
rrGrqdyXQi/rxba4Tvk1Jenkc6hP96HmlKt6T+BH5z2RqXVEzu6GNSn7VaM7y7Lo
KYr2ukv8SnoEJzaKyeFzVU85kzMDr8RC8XdRFK9ucAwVcyiSIPKjSjIn92hqB/GQ
/G8Qsa1hVwx0mNJ95Ss4n+Fadzcw/MRHbsGGx2NN8P/mnvBKm0VCKP907E2u2J76
zxhcboiIpLsSzjmJEHHRZyB3Q98j2Xxiu6JDE4wqcbw4oBf8zz7CN6ePhnfuljB7
TKPFu5U9rya0JvLVY0j2XBUrb5GNTuk92P5VKFNifbj3Uu/dOVqTFJ4XdwvKc61A
TVoFeNKDbKy3+XaEzni/xCLna42+8Kc9tsdUJI9gufNK8vjuP3LlJsAo5xOuhRX5
x/74IHtEg+0zlkwCbQ71gO0z3YynGvWAIGtCDYqbA1uQQx0BRPoUAmQAShkWF9b5
vYVlD/zQwl+3hJpPib6GLiWeRTTi6Ow7wIFCSKp1aR6hWg2o3zGlnIELB79FAYoy
dQ+2uGzHVPm9d5Hxv6665fr6u+QgXUegAke1UCD4+MXvILVKkwazNpdI4KyiORF7
/annXz/pH6U0URM5a2FDf+A0iLlAF/Ralt0+KyZ6k4Ov03lHBqySvLilJ+5XgoCe
IxehiCfKCJoxyTFHhtTimV6merkv2bJmFSuEgOZ/HCyiTQoosbU2bTwybcwL8xWl
BcGj2+RAyrOImStZhQkn0FiIth3V+kjTpAGdCoZ3OxfSJs5R0XtyuSEGxV9qL2HI
hEtnPd2aoBGBec0ML2FbCsHR0yTJ/sDKuj2bcaxrv4g/wYhIJuC/q02Ri6Vu9ion
2mmHGyVyQ5BobzgVZhOJbIO743W/0w+cPyo55y2ggKb5hQDr9PpFvISMI7tgpmZ7
VrKBSDn4besnufj/O5cEUypA65vot+puOGJ/bjJupZ0+qcCZX7KhACiFCoT+TAtC
61rj5peNPQS891vTU6uex1X40W4/8zB3hAZW14bmGupuAA0buaJz82XHMpioFmUc
qsTLFjDXsT5Q5oABl3daK0ROyJV83yKOgOdgi1GaV37WDhe5DfdwdAJpee+c9+FH
UsgWQByRCjdLLgzl2zGLcu1SuE6U4gZhfkO5wM5uBTicnoyyb5ow5gsfESMpRs4+
Htouw+e9HOjbIKTg+lAbaNL+3Fohze0HBiXidH0BTJbZ+GabWU38YRauK2VUHzJW
6Ktv7Sb1HooIdYOWewrsqEchW1w6gdiiHpYU/pAYLtYM0c6tjfYx9a/qUZQer3jT
vXUzAxIIrnQpNjb1+XUAlo3gCxrg+siV96TwouWxpNgOCDrSdfP0YeoswySLV9bE
Ofcyq58byvbimC6Gqh4CDQGgmm56lGLUeW3DnCBYVACIDMn3byucbe4iUPELGPL4
gcFpATBFQOkvGEbLT6TLJlCr4XUyYJ1pqvY8zwLbci+17wjq8cxTDQ+2IOVB5DYu
ZcsLJMD0QBeD5LUxwPq7/qnEWwUH0xumrJp0/9E38wcZsUk9urUFFSswa4HZQXKu
FdMy4a/QUQflm1elp1/CO9v2i85UvfzS7YNVw+PzTtjFhx/KMKhqt+VxATZX7WsW
DYAxQ2N2dnFQnFhyHgAndAT76Xkud7VOkkbbyb35uMI3KMKo5wxVQZXZkXqJ8dwM
TQBXhToCHN0hGeVr2B/o7pyi/Dxi3UDuzwRjq308rGKpd0tBXZna8fpIlyfOyTq3
L6n2TVhT+wCF7l4TbVICM2b6ZAmxvK+zgGPAC5FJ/4aFsWIayyY6vHOS+Y9ktcRb
40Hk94QJD3M9zWViZU+Y4j5sC4R8NtUzmS7u87UfigsR1LJ/nHV1FWeAiqmuV8IG
dNyWs2xi/0x+qkN9UQVA7159oZY31vdrP71Bd+IjU+GsuK8VyirTWb+wgTyF76V3
w0MQIFV/weebIOhJTaMOeXeK7oNM04WdsxIDwkhtqp8Jxs5kLYHwggdrt8R5Q1aO
cLwI/OV72uT75NvuJx/qBmdLAha90KlNYu0mhAn6FIPcRQoOea1PkLdVEho+WDCD
+QbWocyTa1YFMdFUQWmknwdKGHjswevuKaSItay64NyXvVrFKu/8N4E58r/4xXkW
PNd8wgr2GyN4umDIP6pb5ZFhWfCwwmklkRd/8EWA8IOjP5pO0F2BHf6AIbOxAPsa
mozT5JKnGdn5jUcMoiW0fIWZupSebHheHTOnxObGgQTuQDc+UzoXJR006GtKy37J
PhkexEJScq7s46fSouhiu9fMEcA1UN3Iw+8jjw+ApyvDTOHZyOg9fYgdGBczdkkR
Nrgd20HGtgYld4OUMI6+Vy9StK+9eaCvLyYEPcmIuyLcr8qeNesn3ZELGwZr9TKQ
9Wam/0KVtSxqDapwaT+eZOqOzaxtp15JoeIBSLKLUyvkYTZboxOIdTOE8eD1cwRP
7Pc1EWOsC8yRSCVxnSXvzwvPjgAkQamIT/0Rk20HybHxFw+44WqCau+hP5FVXHCF
Cjgz2MnHOQCUXRpPo2M0AO2tfpLWZ866ks+8jNb60r3H2UoMraHupEHLHJTDyWo9
btlcXGzl3vLsEQ8yJogeRYgogC/MdknmwOxb/DFFl6Gat4hK8auNJDjfMxmWTZpL
rkZd9BuKiNtaf41uIqbKkVZDD9hPKZwytDzLrAu3ZH79i7gYI5VXnw38Wgznz9Ko
X5pb20jvxdf4GaylCrmvm8Lad5OCCSDkm/g4b4oEO1n+vWXRd4bQDqlOcxwrTiqb
wPr4xNE23gvdxWUJyyAav+W+ZBnfoPk2IloOElCnLcKt5FnvJFWtmGugBII9Qhoh
L7QhXnTuwEFDEdcHgwAJn/8AiPljbukjSXtIFEv/s0G+VGcIasa9NLndOybR35Ud
QGqT8jcncNe++pUeizzALeZSkjCmOkZANFT0FESYCHJsqmv/prkTQTdX/7auhumG
CHxgun2qfDWlONkqyvpLAmFMDYEq+xFfw43GET6Pms+yEEokqADYapro/2X2ZUoT
hYRIrCrgxbudbloB7OQ4jW/fTlx2ii1Dt/dMuybNxwRQmOBOzpE+e5DbJQQwaUtA
3RSfzzJqhXJMXDwb8c754IAxSkw8+qo5M3lYVfdrde2PL0YdTlgejAWSuK5DP4PI
1XNGOtuByMLOGasgytpvgU5OiPzMKqE0/WBG+2tJEPBWc0XOtpl32d8hKBfO8a9L
HmdiqEct7INiTs0xW3G8hLqx3Q1jGZhDguJmFb88jLh4gFgNYlHhNAknzj+BXZQg
m7o1MXEHUL3c4KFwEPv6nHo2j6BygXgUapNpXu85YYEJzK64NNOvW7jjXknTgZbr
tNzQY2Y11KSS2Deond3Ap37P57UGch5RJJI+rlqpab+k5aj5zh2FelfIkjhqb/77
DOIXXncEXNVc+OlwsFFvr/VIlL5pCJbB1AsLgLbQgGWkm+3xilG+N4Kz6Da4IA1w
eb6BxInUHrwq71LrqJhostxt57oDTvBC4Zrk9ZJlAqG+JTM3aB4XWs/dRQlnuoiE
axu47ILOIT1gyryaLsSNkKQtIabU1oeosgSFtnQ2iOCYiL1vjET23Xn80UXX5rn2
KONxiX20uF1DC5GDUmHncS3CpWe+ap13Pj4h5bbBusVOqkY2cUScan0vJWswABoi
jpcLnkHtOD+fkuqRP3tYFbjSFVu+gof8EQOSN5gVn3LJvolnQWEfZUgilsX033Qo
gIeigRMC+lVLfj/r2MNkZAo/QdGsbAELwsI+BIw1v2R6AR5VA00B0mQyZf6yKCvy
2VNIREsoexfELZD/1ju1yVXTa1TYbiIJWHeLRViVnXSbwH5Tkmb5mFWmTqUc3qqT
0EyArdTuhYIq7m+H6AKkVqBAEP6keZ3EhW+oyOnhENawjeBtACBWWVxVikPlTYWH
f737S1tCa9E8nGqBgSqMgveRw465f2/QnsqCj9cPjMYu95ciRUehS4nociOzdMs+
uAsaqVmWhApodw/VZNuBLul7nVmDDMvqpq13EwAsJdUIMOE9vjjUsy6SNNgKvaZS
XCsVUi1PvymteNwMHgwV8OokdYaH5RYjqc+oneqMJmBdVmGRukVM8l/vT40EnL6f
OISG+xMIjQ7K8hWvBtF42CLMWhXNEsq3Vz6L6Wl34CupbgmXwSC6lv0yPSmE0y4k
dIjiUf54eECsUKJXzl5G71oc3qyijztXpIGjLeeCprARAjwCxpBL+vGXcwy2xmzk
XTpTLG7ASF/sPw8EgiRWs+dcVG6KrSA7ljcvbiB1LLle3DfSecXynaWEKtiqIdQm
tNhaw/K4U0IaBsEFeWvNGjGcAbkN+qJ8EUe34pIZSAXyv8B0F9yuKNm2GF1CrHkj
ltsKql+mj68M0GPn5Xx5Lg0Wzo/M/smso/4Ies91RDYTFhime/gD8XsySYduPP/O
5AhNkcPBHcmvKO2tOGiOOradIAWDq+tgPMYmpqqYMNpGW3BeOe7j0PFCv8BSNRu/
kLe/DucdGkfhKab19HZzzBKJI7SyEIbXqHE7L4dgTT/nCrsPGI6jhIs4PpBbGcnK
LBIOh6rzmZbX8pHvno9JzUryMd8TJkWAg6KUbttrS86fGt+aVVAa2YrgaukhHJar
cPdo0FAeKPSafwoMYXv7EOqN5xMsY08phtEOBzSvOw/NRrgCMyFuqrb6As4anmqu
4+SVn9pKkJH5OjvYJp19hdNy/+oU7YRd9ncz0u1iySMW2V4l43kqz4flHDsc3ttT
0S7y9FtbobfnXsVcElvntxZOYqnPW/7DjJrF8MPAXQwd9YlkCikh8DqrWWT+kqFy
FZRPPKCLlB0+TAamIIsoc/y4hdUmlVn6T6We+sp80SvDZvMeZyOznLmTYbDfShZp
IcHdpKfGUDeJm+KkTevOCiA68y4z2idrLQkTmJsaorjOuRcIHnTj5mTSXckfEWfr
26j/ZG5TuJiLuYCHq06DpcNQXcfHwrEh/ErEf8d9/Fi0XDcC+WTG93g+oelm/wzR
WTuposCoYY8f0R8fGVlc/TqM7aLWKilsgJrsvoUU9Z0DyPjpMUeQRAq+jIUZCbu+
bQE4KSCWIt+MJINTnzAjCIuFlmfrWW0gGjF5XZ8DcDP9lJo9ixUoMBUzsnZgnNy0
c3cJbYJgwCXYzJ44cOG2PtOEyznVbIpK60otVoRpOk/601j7sfdd+z6n/Pv3L8Sl
6KTLBDB88Eu2r36Yr4RP/EqOcSWIqoqMIHWCPWREqdCKc3O9io1AZSx3PEdLzvTX
nnX5OnPSAiH/CPnY1NGCB3P/3dns/Qbn/UtIfY9KdEguf2Xi9tN4foOpeWGOjq66
OP++rC7dZ9zO0ClqBuaUzDJYFTRTliwx/DNdrFu/3VfybDtyZHnJG7Uo3O+KqiKV
KWWmMgK0ReEZiW1kPrTXwCXrhz4BePLlumAlMGM8tS0VO3V0LWCe6q7pqKQlwDyX
5/RNCZSPRGuNslUT5GYdOkPOaPt2EsIW8kgTV6JOux5alEOZuOsswW7dDAUMrBT6
s6N8xXOwSVk+qVMRGTbEF1uKek0Lrf9opIlyO48da1n2VEpOaVXFG9BDMMzhZ4AS
y6zNuXgNSu8jDBOHGJLh7F0C8Wvcgq7rAHacIHERJM02P6h4ixbhmvdJOZEyvS35
FEmbNhOZuWu8ZIM1pqZWh+ViG5RxGNxpkKJIx3ES8RaluOMSu+hIdapyyvKweq3A
9Rs43Ol5LIB3DBJNVTDEhdrVguCblT6jEciULpnT0pFCSkYHSn30Oa4ShaXUhFWg
wddOoSDQXHh/i0RfVojL5UNMQNx/WRDule+RvZzHZruM6sBA6Ytqx59Q1tHv9cyk
ladneJV0fsxzPxIHF25Jmd3ahy8fhsEtawKrzSUTGaMKV8Myxm+GptrWWSzZQU27
y4SODGYnN/OFiNa+bTogOo4AT8StnG9t9pPBloIfFrPPN2ucDG0SMJju0jWCLn73
ikJgnpemcEc7YsX1zYQnEHiXOB+RdpFtnxU6/lkZ4SkgjaM+ADjIcOEb9pIBUZ1i
yf45yQ8lKpo2KiPFcIP5MXX5WKT+tz/1Jy1qnDXAez0K2EqWaST7IcfnG8KIe23Y
KFTcnSlVRe2hb8RLsOeGf570UBOAVzLPR37/CrEBNhh8iSfEhT9ya68bqvqwNof+
bmS7kFSKcYSoEvpQxBGFdP9hA2qsewnKwtZM8glApTtIMgmdBuLGV7y+Fc722DSE
M7sD4fuoaPPnEPpdGHAer+ZBg0CmU/2S2PD9GLrS4PumsKzIloCzic6DsUDq86J5
WrTs0xnb2WMZr2mgMckBR9dwLXC+gG76etuTfMPvU08T0FnL3fOF5xRh4VJ17gTA
tP5NAnkzYKViRcCXkg90p+ANvZAdFloDl4Z/BgpzaNpJpjvpzCjTFrcYv7PXwLo5
UBBrPP2W2X2t5ReFfPFetvAB4I0APJPnwqAS151UPPnv7jA/mrzpTrreRPGf3ZoN
u9NW3AmYAB1qca46RmQO1PQ9yE5JFKazT4HDRiLZJfnxIWQEywXDAPd+IZWJCf/H
jsin5C1qvUfsjx7QTTcfYn890wKWjijvSj8wxoH0qWzpJuefcbcOtA7Me6+JCuvJ
whukOK+RgPePUYkjIYJAmOu2vumBTPA4YEFWB72QD/kLCGS6bvjZxAirvOQg44EB
7batmL28pblHKtK0KPCBenHK8V5CmBCp6j3LPCLvcJINeezULhJw34v9ZN0X6zKA
LBoBw88a1dJCZQ/fzxFpghnuIXaKg0a+4wV7sUhIynHlMPZdzoNNqWM2zVJEHch1
ZtuyQkMteaPVWBnkmBn3bQHBFPSiu2cjflTb48T1wKon4mB4eiOWB+3k/41YtQab
SqN4aejG2KjeQJ/WiFW/ifvfMMhWZW7mXxmcHj/GbnoaZVTr8YtsLmEzGRq53Iki
mbyPlBuU849pMYcUKo+0OernhXLp4wH6BRnmcRX1OOF1gQEYhOCEoMtDSwAh2ZU5
AhVljFBCbH/wjc6OW1IFE2V3U+VYu9B+D8k86RubHpPIKxMfXtxc8vtd6jsOnnFb
L1L828dhM3BL4WsGthDz6djDkpES47fRJK/E8VRMDE+XUcRH/m3YchWJRsVAK76C
ITbpQYUoLbtSg6DSPFAAZb7in8sRTiBAoIVW/+zOqixE3HK4bqs3VQgje3Me799v
o8iipRbTSSlN422WKBSeOS1rTR31vuNm9SN076RVBHYYIxBHqTD2epCX7ZXfxj2m
ui5LYsL+uAslqAlCk7geCsau+/92UvrPEi82FeDf5A/h1SUiLbkd+/Xch9V+7KBy
ZdMysDybHImT/IVNz4Pxklo+YygcXA5Jp348qUW5X52fBy5D6cZm/a2TZMha0mP3
YGxC0UPQWCNKudV5g6aPsjDqs7WGGPoYe6zfGq5ABw4eCdvsOVxIkJIiE78PVx3j
cPeZkwGZmrvj/c/eLM+pd84yuYtok185PdO6UIPq42hJzSPyNPpudRn8WezebZHn
Rf1ihvLDOndzqvv3VR8orJqmwZDSmgJC5+rQQnrwFMCam/RWGH9VlrO4XRE9U+Cp
NLyr9kV2gJH/O0TJY1ZpWF3UW8ygVA7A794Z+aUdpY0QUfWH+MVOTn3ISAyWgukJ
WesE2zkOBQlw5J2jf7R+wUaKLHAc+7REjSe6dMbNvTixK2LxThNTOsy1RNsKteR7
XZoWQg/qdIcN1zMITkRXFWX+bAmHTcDy/L3QmFKEbArIEodehEsKRB+ZuWBYu1U9
IbEPxmWGf2+tGW4rNNrmM/CrwTBKnwFpjYPeGw/xOR2HGfrOrAnMCXMdfDrQR34F
R85cP68wG8WZk6u/vt3QzWLLwwMuJDrv4wNbJFMv3OY5Zy8+G+6qHWo2IQoET0KC
I9VMjdcQuuRwexhy8/h8bM5taAOICwm6BmpmUheKyjXaSYz0NfwLGgzWh0cFeym6
lNRcTO0UoLP2tXtLFWjNEx2YG80j0zs0ZSZ4ZiINxWcKEF5aOoX+jVfO36cQffau
Eosk6A0ZOUHsRhVOoFvSelEswajfkOqxQHUkBlbjY632IIJ27zQOrFr0VM2S17Tj
irK8uieyzLz1duUpKBoQXaii6p4XAv/K4OBHbkl3yU22OXT9+bbAQpG99KV3/d69
VDkEnUbmPFsmO+AIO3ZYvL1PqJmVRKlJl5D6inIJJwEaY2IvZ/WI4rI3wminlqc7
m5MGzd0JlwNep27vsz8H9oTx7wktnub4nDfoa92v7MF3lDBJmUMsMakJEXDd9jns
CtqPP3AZ6kZr5qtStf9qhduRaCiFC1jB5AP8aIosa8PK1jz0q6pK3IB9t/Oq1MQi
AzjWkW7SBFXYRNdQFuALT34jmA37WvYiINQ4VHIYupfFJjCUbliQWls5SuQHTtGT
6n1CRAed8IESsAh88vu0XFxK2y+O2kjB9i6n7t/+OE/yzM8CR32ZiDw8XD+NU6fl
6mqJgi1YNxrrsTdb6uPCW1WoYJ9rxcBpNB2xxVLBH4xBkgEZrHZmgt/YN5184U23
ysYIPFvmck5ehyWt9ou0UFNNkOpNQ7XRg+hpydncrypm7e3DSWhXgXYTYpscEXo2
0sn/dbPsB2cxoUCFqPMDJ0IaW/l67UM3ZrW/LzUobuuBqETdsZK8ihzl4foEn/Xe
exOZNVeDdwSZo4aX/bIZL/NtO5XOHeJKuhqA6dh3yda9ssCNyTDYmKercL5at7nV
4AtvqhHHFnTB1rIAsIZ9ZUrcto/2zW8OIhNe+BAlXVxzz/7v2zBjroc70Tw+t53H
WnztI6orl+Gl4GQOeYpG/cPpt/tvW5v70vIqAujGbv1xQRHmuMFBoqyjisSaPuo3
xlE7pEF9zSMWz+wXTtyOchmhV/DufhIa1bPk4+ofvRt6fNNWuVHLJA3yuZbFDiP6
QA+NKhliFkD+Hr0N3zw4o+ocjI5aBicXjscih3eEshD1HNEIDRj2mLbjXu7Np9PW
jqde4nypEvM5XF+IzGPb90g5rkX/qPxc0jGDJq5jCM9fVkJOKodpa52LUskpiPOX
ncfR8MT/+1Az/8vDwoTTrGVMsw3ratuAxR3NGCySRoTg3YoALM/nTntn7HmrxHSq
e5OCrzV6d8Cnte03hAhUL2C3XCnu+oSrAeA31Llc1k1thbnISfz9A5A1CQY+XVgy
Qkvai/8ZATna7IvufcxkFh8aGvWfrmHEG4JE5HE91RBxvQ7JWo/o2rG0Y6pP+kGG
jNZsBdQ/XeV6YEQHvMRBslSZAxmYXHLeT/j2zRKb1fioemNaVTzrWGD05hxV2xJX
0shb/6+Non92kBw3GrfXRKEICDI+oKQyCqd1TLNx7NpB+aNGd7DbyAP8a+rJxZg4
O8ADju3CuTdsdikTYYDcdaXnE8ZTT+Z7xR1zQn6duNYXDVeP9dhknIFycYkg/ip3
NLDiVJ/PWcZWgubt9Gfu246KiWaXZ400+n/nyQSe55pPcnSRCxiZlUY6MtqYVLGZ
c1gokuk7RyQF7A8pD7H3hCIsLy1r0g3ICGh5RLsy/KohWtbYF3+eWf9Cu+rSGyMX
8jWjkoay+n7yb/IvTfql5ii/tIV/2xGuMJwLgFRDA7qMZ/2Th0LPXFo1IPTcXVDd
PBH2+jQZPXlgORjDOT0H3X/fxvW7qxjpHqHdMjJAHpwldRaGGMDF/RJJuLsm6eWk
AV7sdMzkkOZE/RuDHnpXqK/o7Vpo0mbhu+19aFFY0Dej3XwWkY4+P+9SaQ5E+fIE
fzk4e4+k+70DuvRbev790RRMrslvyKnS9QTwIgcBmhZA1Xa1y9mjFglP3OT4i3is
dGGoT0BpLy0Ul6qLsHPFXedNbCv8D16B96Aaoy5zHa6MSlGnLvCkwpVNLnqn9fP4
dhLHT/GnBqgAzdSNr6cuGRLpo3/ZOkoGf/1okFkCicz6iH4+dPFp3oXaZRNOHWNz
nDWrAK6HLhBTGXcZQQpf8igwnXbKWexuVlevNM8qxygeJELiz1VZkqYfDo9Mq5RF
Mi80UOAC2lM5DWJCm9fumkl5QJvtgoG0MqaR2HPgvrqECaKauJts/R3lmjcPdpW5
DYc6akmGKUJRLrJYCwlal6xD89pIHCP/ROp3fa3tvZlxjlAgjFw8lZePmhtDgAlz
AM4dNx1c9yatuEMpaFTeiGLS8NF0VZaeedkss6GR68DGnCMd/EOKgEc8l8pIMTw2
JkORgN1CHnGXcVU3k9AWzalYZzWGJZSt8YW/Dz/5/qBUOaFVr5xnCTmrDmcTh0eX
8qZIwyyZVTfZBAlW1s0xA8+kRIMUFFrzqFcFYsBX2rpotuGwALtLbcLrsmHSHRe3
jY0KF+hYvbRJ6/L1XrsHI2UWHldQaNfbfFIQWYU8vvh/lQvFsHxO2df9jXyfY1n2
OEhR3pdgZniMl2TPiyQswCU3C4aZcP7q9Gb5TxpEaiaU83VMd3mF4VNmphUKUmx2
cRZS4i3xL9CygvWD6TVXV6HuF/pght+hIqA0wN93gnaaKhnI/0ZgrsRLiQe6WpY/
CGedg/tsNluFOoM+gFz85fLhkBdAyHGLDzLABn+MVOANGCnT+kX577dGXzIaMjyM
UqhYAxhkKXsUdvwU9fvd9OhXaTUl/6DU97NsWDp1CGiYVJdNJEy0yob+pyKiTQFn
EBgcDip41G55Wwix4bmsF+ISOfn83jh5uKvR7S1HBj/1GA2WatfbMrNAjSojDIa5
lH7aUFYlnNG8jeI2yFMBy5Kp7VQyVZCSLEVtnCbtOuwnR0p17xOAumlQDy1AJ7+V
`pragma protect end_protected
