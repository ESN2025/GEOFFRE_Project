// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
m3zSrIUVMfDO8/4qmPI1vX/7pjF8uTUqNbEevgjcYqfI9FJ6VBJwAfHyd1tL3epn9sNaT8nYt5ON
sHcRK+GPHpOyNpfZpFCjiJNwWtjbL1rxLBhDb57dHz2fLhppzdidL6V5auiCV77JZ4zgss45tIIt
9N8rhcee2p89BgKcToLnkoS0eoa7vwSAerbwKe8RbLX3DsPe1AZyy2CKeniMYjLpU+hpZK5ky+Ka
ayq5E/VTWGMPsdSCRT607kaaOI3qjwuZEnFNzSMtVoNZOPNpTGDcD1G/UjnFGCY1XHno2AtWEDee
/i3qrjGJAZIFrKQqXcdZeVsboGV7FcKemjcnMg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 36048)
ulM9xx8othJKjUe9mU2nk6MNfPkCpE6VotaVCrCqD33EkYwC+ATg6Hs4dvvM0n9tm8McVFs26Ek8
pn6a1wco0/84VRZdalXjPJbC1+uIyUIYPLR1mxaHSQ+QZ1JHnee3YvKvV0Iz4h7NAgrQv4pIP7up
Tu0+sdEkTheKZO5YmOz07ms1yJDxuewq2DhX7qUi7kwQgq4kCLNe956mfmi/p0rJtB1EFFlh5DGy
K0mckpykmsBBhUBFePDpE81XkdUaagr1gXOI9EUwqu6/VzpXI5C+fV2YhCsvk2TRQtyror0H0k7p
rbm7nrGLMeJCGL5imTfkQwW80sLXUaPjXPBKOMT6dNLX2WLOaFIIDTh7y/0gVW1Br9L4OpuP6p7V
CeRtEaQO0mBXaEfmCbpSGuZsBzuUpsx6sMoAvpOEt4WVHt0KJnWhtqp79y9lNbLufbXWyM9uKveL
eVFurRKY/ZV47+2keuEYiiBPfWfQ2dKyyEbHBHbd2/7NTsGwTDu8z8/cQFbTNZm7A33zzOdQhNYT
ze6MXIOxm7vIkw7hWO93VOpeG1mJUqBBDzCl7qH3SmHt7TrP5RtRTJ3jDOx7fiZZptfz2zdGYR3l
9mswBNTvi8QZq5vESNjYShCq/lk2icb17BSjyqN4o/cB6cDhr7ceXfbWOuW5pQJYRLUxpuKQLdyd
fdwPZ7CZjqGyjqG0wA9y92jMJ/SNmhaNUoR3tISd1bFhDdEoG9XNNhY+8WNw+G2ajXiRbOusk6jU
l8xLlQK44FBNzzCXlzadoXJ4NTttD1ROIhXhnTy5dF1bAFVgEwKlx3utNpzN+Frgpvt6KS4VeLcZ
rxLqSJk5rZw9yXW8BbLhrzsNKtR4nkRFHUkGfNmGT4WW7gq1jhANrbKSWUu9KuOZVv57K/97A82d
PhBtkr3LZkX/0QvIqU5M4H1TBt2SXgc2BH/Qgs70ZVEzM6aVM6bFSJVZSsfy0XlPrO5QdNmDMsKZ
N78eX4tRaloscUkklXhIY2o/t4rYOwTWwMZunwT0IXaxhf9l6QmdJ+d8QTvuAqnq8ULD8SglJlkR
haVcx/GRoi41puQg+vJu5tFKikA9Xtnj1KSWCV8RpXDvEroOdZ7eVMmC+krOzEe6VwkM2reKSQ82
O9XDUzzUQJwlgu0AVQCy+QRESYwKAJwC07ddjawxyAsT4Rf9ITGw50Iv8aYt+uTmq3FXq6HEfUf4
OgiyX8aaaAUbrYym6hr9meWO16bwBfawOZjb2GSwnM5j3opgE/kQSCAJTzeBgVxDLglrwq2UkEbV
fBmRDue9hpDJ0Doa0HqGjSVVoAalM4vaIhzD8xnBzTcfVOVT/k6V5O5cPWddBHJIUrgUpaT9/qkf
zD/4adpndc8is94K8ldnNzZckIl6WIjcwljRHnlkkg6IJd7ZfX053oC1EJB4anqpPxzyvsqZIBc6
VzABfWcOVA/F9ehzH17veV18z2DEkAlUATbIEghOApg81GMm6QZNPAA8myMZzLDus+JEc4Z70p10
hO5f4fANIsPEkorf3MjhslLYuMk+mNGVHxhXkOirpRYdkItUCsn2sSktSUIvK9S1OPuCFwA5cHad
DrBQE95Pge3QDmgjvq3fv4/kayp6aZrBvylyNkHlLHg48I/Ms2TAWTyqGvOCRYPLm+eQA68fx0xt
Z0D8QKj7qDfFaz90Bj42Izz9Na4oS2nF2gNfDACmhwSVPVr8mbBg2ahZe33Kjc5g8s7w4bX9JVj8
4q8qpp23cmeuhPfIWU1az1JIncpquR6/WbNFTzx4V1fNvspcTtvEGnjI3QtTowwOv/8y/k8OEAYw
ugP4Jd9cCyfOCy2jj8rKm33mFqBZgzUg2jEBjw5Z2CG4WD5ev85sTdRwvwydsVulxxJs93AIHGjF
Eb3JEHJiw35Xmgu/xJ7b7VMN9lALIRu8UDhs1gjgpns7w7eUeb1K1KpMp9FFymEl2Wh6m3OQOpEl
AUwqONWuvs3d/qeih/WaqAntKpgkgeolH9jzgW5SkaTC8Foy5uenyRq7k3ljwykKf44JBmZhGq6D
lSKzDU1TwfPRAX6+qtf5pNAHCYAPLs7AjFqprN0UztFgOfWroR47YFCtAcUC4MvvzIidzSSCizxc
6HYwq3PseOEMln9rCuz/6x6AG4Ksx1wTD4w+NuhA12S5t+hldcxCwg2aXdA4Ac/YT3cOtOhLgg8m
cTjLpcgpkvY5dtdv1reQDLXbO4cn0o0Ta36kGOkaskXCFeM5BpnBFdsO17LWlTqJRokQSg/OEeeF
QsCvDOv3xFNhW9zdsVYUnaXEoB5aozkedyDeM1IWwcIawF2TGekKWkp6Ck6amOMuLHKxcA5PY5RD
WOAGMyTDTYw8aBcyUXSAitsl4GB+oUOghk4ErH5JhgJnSBXxZcZBax2pjL+LviHyqGi9FlU3pKyf
1wtEQ4/anKuOXVYZCdmfdRpsNEQpRlnZBCHR5DQJhU5UCJ5DYgmwePPx8P77UagGW9h+XfK7J8bD
pHQlDrcLRfKCYxYlXCp0PbT1iGApGx6fJK096CXUcnx3I/ajGIN7HDJEZV+30JuN2KP5AOCn2iSA
BQKIeGe+upgiD892yfrdpuX1+jIuYKUacJmaq1On1BIpOUuUmKtkcrqY8tD8wIWuHoF+7FfLag1A
hVcRIfwBjSPrITdPVxTFWyQwbfBtkUpqbR0uUq087UyMyMl1bERw08HB4wSjGiiXAnjXKZk3d5w8
Sn4r73UYaDK2ZLLwL0BvwheFwFvtjNTnR8oO076Jw+Mj3a5UIgz0KXpvZHPP5yd18/AGYhFTZV+R
2gxWJLSlKnmx3MajAT1U8TMeajlxNchi1cIKOIljOZpnIIFMuGv7fPA2sJJX1ec81WrETIHHoPx3
EcqaTmEjLRvOM1sfbNPU/vcNmrAwSjqR1yk8h5hlREgOfBsDHb4s9keOAPHQrXzxcJNEcZHcZJr5
1egGwCNh++RyZGNmuXiK4dgD+NFF8N0t7N0ftsURuRhV3CcSkiiXUwzUu0GsQypES26fKln1o6L1
RodjWQr83lBxSFRLK7htTxk34BydhWzHfX2sD11R3dgH0++CPJfZOyDQ3Z91BzrowwmurLhlyGxK
Q33fkrHx1KQ9XL7riNNhkmFiHpPjMkjuWR8TbjbvicpCurduGFwIcj0I2uRHBfDggbqtcI/CQ7/u
ifqSs/PA25ixSr0j6v/qeewvxtMfn27+34fY3IQMJ06j3bSyoARUBVOwBXdLCTKGfVNZAgYzhm8m
F84YtgtF3Fu6Gn1P4RElsJPl+FUjSJ99IKW4m7dGyY5DE34qzKSxLcunpyyCVHHJ9fdEwqXAqEr4
4TeTNQpc/gLwSMwdsmOlurofGyZs5iKi3QKcMJBrQvS0PoUxhR3538X/3KIlrlITnBK92CKNyDL2
ITNS2NZCQSbLfvl565eyutgCZ9zX9lnI/O9w4uzpqY/FCZTB1vq9fiNBBzyDd1PTQspiQ/YZyfa4
AnZgzJY2W554CFlrV8cM9WCk+yusQmv5sqmtKH2PBtpMfnSISXA5gUgUkHtp5Z9+e76mQ12QKh8F
UZD0IKVYCRXG1DSxoj3wYhZEMbK4lcyvmUICdXSOzLfMnNrORbln+FOtfxaVt+ywkPjD3w5AZ0jc
XFFQjxcDXQjPsNzbVplgR04F5Uswnhg2PFO1UF/LbSnFoH7nz9r3jxW29OzHSwi6GPpIKTxDnO2s
XX+oNNPpxn2oI5DA+CLXF8BcB65YM376ZRFRGJMeRw544b9AHeuAIXCm8Gikn4J434XpTZlW4oPc
p4A+TOum43YPvqz3bg1QsNujm9tvi78C2rT+XoO1Rx9u/2TIQycMROX2b3dNr+p32GMuJtPbTKHt
YcBTSFEdPp0x4CIM5++TL3ERFUuvbxIpVu0erfSpKuGKtK4QrkkxiSVrgkhRTD/67JhZyNRT9bon
Oo8tP5acyS7LYiSTasxvpR68utmtb85nsHd6P+vHGIz4gA4W/2PlQuZk8FH7DFQEJTiTCnm8LY5u
UMTl+Ve8RZzuTgWchuVKQynyPWWoYtF9py+iVwBrmUzg0YMib+kPErjv7+c62dYYyEMyUeUnnnN1
fn0BdCDeLM78HCtWDc4xAwLv2wiMYwNqSjwqBx7F2scwTKiJXzygTcyL2hr+hb2Hjl+AL3qbejq3
mchdgqSbfLCaZkKGVAxEwnkD/2+99sz1bH7h++0XhynJLr99yY1CZ/yD+5PVxjbJESC00o6O8N7g
mak5k6G0E/qQTM+erS4zvd1WMqz/027Xu+7WPiaEMMYcoAmBKLKe40qFpSMBDeli32XkSfTbNUWu
AXlLyCcg/BjWVoTvMzAeUblFtoJjCevhJkzvV6xLPNuIRHtrl8aVfS//A4exWL4S0Ev6ESXtjaFw
062HH6Vn9+GELPH2//4Y6hHTtg0IPn4TcYeuzpGTcDFIed8yj9qIhFJR4IPtRxaldjMu32H+6eaC
2V3pP+A/48Z4n7qVR+wslfSO65ao/GSIzfOfAW4kyCDcTV522/P6L5fuLZUnr3LdYorWYbCutJ6N
7moZHCmkLaJYTOq0krIIA9XKdguN+wexLihKy3ot8ZWRGg+q5t5Ls66V2wRWSnX/5fogYbwd2diL
jfpHqv2jUhhiUalFR2XJ0UQIQ/16eYpicS9tw4T/TneT/gL0hBiQQNKmEwQ4VNVpFVN51oZDm5U3
S4KXll18b1nTteV1MQn96kucO2uOqO2fwS2lfdzVd/Y4grZRMGSEb3wy6dDjoDtHvYv8aebXQ7Ca
V52QRHiUVE1CUqlYi8LU5rMAjj0/BRgnLyVUFMSZRNGsMkqyLR7PJW6i0wsXvuKJpl3EQt1ylayX
qUVEljdJFJv7tg7Sdjm+rbUEt5BJ6PVf2yneeZImDf3ONYXKY3CJpqX7vRUw7b7PaAdP5DboX9Kh
tbtKlavHQdXJawfTASN2UxKyymnmsFvVDb0nxl+qOmuCABfCXVaRrQj/ONbJR4GGu6PDwCURA4NV
Le96EfkURUpeRe0Yo5535THszpmuAYes+t+m6TfekXaU8pNza9gyGA0Ye8HAkZM+v0uJyxEV1lhx
65lVsoNO5nY072FUHwOghe6TUoH3whdxh5LC/Wtgs+0P60bxfi+gPcZDr/5yWZz1LPvHnSSfSoLF
IZWUcj1KxzDW4pcRXNsQHdJJVudQyNAtWS/cOzXJKRItpg5DCYIrtGV+nzTMLZCbmR96DJOD7WT7
bjHmD6RvujPJY9WtA2JuS095NYJ+rrIROET9RN/+5t86o3kJ7LMnK8Xf2bbVdjizSTFoiI9w6wYs
FMgWSkXtylmstOdTOZ2rrCZBvJz0eN29IVBz8WzOaNO4RyGQXDP3r0fvl9MfwwHAqn9uA2RNK/bU
xbjM17EJr6eC7ChV+t9v85XcHaWvSFngimkOe2nong5XscPh0dMA034A0XdLelye79VklduVNUYE
Q2S0UYCM87cWTOKuTmOIhMUIrh3rocIudsHLUvUhPziA9VKlGD3kYrrE4VLks8I5MGc6uj6tGrlB
usGS7lhMkIcTiRPi5HEtBnvBNNrhiihzRXAhqqv3X85lUf4ujO64PyAlV5/P6XmCR97OgUTx9in/
tvyRuOmgPBw52stENap8QdmVGQ/PHPpxeKtVvLIp1dPQFRP5ma78fzOzUqFsn8EG9jsTF9DKDmif
zyhhNln3HByo7UE6EO3zaMB4IDRevpSzI9gEJ4E6Iso0RQFJIVOZ1MP9IXwg1jrWJ1R/PVtbEC2L
oRzpdE0QWigTE4A4c2JWKlzaBEc9ThvDU9dqOgfaZGfF8KYucOm9t2KuaSNaUoGwGQL9kqx2SsHQ
m3k2NwCqkVSVXHaMxdTwn9hBybayUkYZMOf9+PRnB7qxHYZOh4eVXTlgZbRobf6LVI/9JyJWWIzP
gi92ZJRBj/6Aw9ewmK5KcaqSx5hmuwFmBy42Px4EhUPyKO0QJTrEPSBn3cYaHDvEG3nCGbvZE7TJ
Sm7zOcM4Ad+oErTyU8qwlgs7hENx5eYzqPKF/xq52nXHn4viFDG85XIzdjfRO0vLf5OMP9SlLbRD
35brZtcZw+hHsJ7qW6JVZgqr29Ce4VE/KfboECdPt8B9H7++f9n7oIpobmS58Q5Y1IgR7QKenz5Z
yufd4vuTYb4qwwq0DCW1XLpCwdXs1a9FazYP+5vyNU2nEme6bWlN1MVPu61u6jadUV1ozzWJ/Fax
/jPQCB+su8+KRs7uHsPwbON2H0bfADEajdCm5z5XIZXjdKtWNtKb/Q7d1wKmSje5Lsp27j0CKhSh
VoUc8wxdffBIFtLubQ9GFeB5Qnwc+qE+G7SDMbGB/Idx8wyEZ1Rg+yxDTd5NFGOEbdM0rm3DYtUW
JQ0LDPupThTGqHCG7yUs5z0tiDjnVvAIist1WfPGmWaEd5qUvNK67Mg2nwkurUTjSiulwOrAIvZO
T3uTUWs8X3yntvTiiGpW48Y+ikvItLRpEatZ6dF43E1wQW+nBl3KFj7IY1mcdB1o2cMCZc889qUZ
D0HEDIvBW7ZGgmX/qz89FCv5Ny2aH9auoDq3WG9+/YnSW5PURHNmg3NSIBFzidLZj31mn8y9hyQe
sVSO6VOyqSMcI5rwkUJohCCC8gCkhmyXO5LO88lG2mkiVUa4OUcmrM4F5jFNtEyYelKwki2ALuQ5
b03iup/a+jSCD0ErIwpA4Ps5Gw98Nrh1OfCYe3rmzg1k/oIksJZKakS0rC/9x42c8NqZl3Zegq8C
wyQifY+6FtEbnrNWHwjYPJJPBIfWXxVAHtNrnrMnqwNNRDuAI2ZeTknSq4rCvUibUCjjJjgwv9iM
82cyOuAMwsmgfhg/3fw07vlfkOBQ9U9eYRp0jFQrpyXUEYdG2yCSoPUWvh6s4r7HZvEJ53S6UTS6
+UcL/YNieJxQOyF4+FmFhstDJWj/jB+Ejhejx8O6KWo59EwuazfEicPnPrwW4WzgHIF7JG3MGjZT
+30kndwk8yqMpn+Z7d+EgB7KL6ANhY5n2A75onUefGGFY+6l/0Nk2wG2nz9V6qZj+cmocm6agDpG
Brqt6lpSJJuG1vzUQB1uAEr5c3P+T70Rwz7hc8STRXWIJFXcVvJtf58fsov8lz3OKypvW8MoFJ0E
hgIVZbMf8tc+J/eE3BNbGRqyK5miJX+4TukkOrbqkaaxDFsUKe18B38OIXNO9G8QrvBNho8QyTCA
hNML2M7+ugQ7x3J6R56DMX86A/5pImMGP14Y0KsCWjAG7rqVzica/olCrqgnqGuHmAhjhkh3eeAY
yBchWmgr9PzpkzE0oPlDdXKybfqyyj8t8wQivChFZnq4Y0qx9ZIXik3IvcvrHA3aZgM1MGZN709/
HhCU01IRqwqOlrQq37CgRgqfKI2t+BvXWSiR6baGVQi3zx0R1ETCfQW3vKmwmDaTefBIr/Bzp3jq
IkFK3kTerbxRtt3YBuo1qaDLQM8nsw5GsALjyx1j3zQhl0xrjHoVhucY0xLnc5uXHv/vlZ961moq
6/jNrogxnasEJSvFNX0aZ8R5eJBNzXnUkZ+WI2G1T8xCUBFsM1zW+EjnwSJTZpReDBX/HHQSSAdE
Prrz0ck/zGS+jSDLLZC0RdQo4NrhqgyZmKaYM35CZM9SP3qJ8ZOXkELK23iZVqG43oqXk/zwaRVZ
0KZXXbytgJLo6kRaJD34nO6VpQ3FtI/BBwv3n8SWF8obHsHcgtv048Op3yiI9Qauw9KEgDgly78o
C5I/uhITeqcHYJPkISCfTvtPuqTHSDuBHmSplcmSjfrTNmmpG8FxgoaraWbgeyaaviKwcL5w2ME/
wx3CTUjjAIp7JxxOj9sURZO6M6okTV7NaOlF2X1zr2eaSp99QnHNSSJRggb96dZExEhdac0Y/qw7
hGTovasN5X1oLPGRSlGUjN26al/LS9Wm8UrcmjOCseTaSXCupiOpHtiDdVqfHeHaW8GfzOCA0f/G
FUx7pgrEDDiRRzkAvRuvtOThgG/ENoPefg05vptpGnhq76QJC3mcJ6naOg7gFGORLHfg3IVUHjAq
bZ0PV3jl7Qwa5/xgdy++ORCAUJ82JYTdAd0f8zvKK8b4z+RbYxs0lOGnVxml0CdK82sXhstIy1ro
6U8SVkapo0oGP+oQF2pRLn/YMkFoc/5BMwSuAe0qpAW+3eCwO/dDoHxQEnwCoEfPU/6uylrQlwXA
Q1dVSW/Ge938S6B6Wn98AHkyZRPI3SImU55A1w4Y+3kAa1HQFJ6MkVK9b7wivxf4hOpax4+DE2ac
13Fh5C+8S4Pd14Jdhz7OLDIat85KlbjBM/DuVJhjEQ3EJvzvvE0DgB/2s6zVa4WybKrXuFy87ItO
Z0o6eoa46YYUInZv0Klt6XKVjEZ+lFsU5unyA5I8Pr82er20lQZ+E7Si97ZlhQ2IKmR5ilpz7P+u
oH8ZDsDEd0e6B9MOVCjErRLK/nsyCCJk1+dGwv+IrpPug/CioXLbhfcLEouyZUteFDZ5uQ3IyRD2
SzKIxHHxvX/W9MQa4Uaa2WjYFyg5PNFQYFeUsd8adrHeGlgY+IfYTyjN7yD4Rv5LiglTUP8wkeuS
s2aMUtQNlR7cSMXOPGd82UqBLIXGAbGvkk6RUmsSk224672trNNEwAYcoE+kJhtHtf5YWUarcILW
aPUghrMiUcYKqnkNWIIe/jNr0seHnrgmXTSIfy27f/mxLOC2FSLrDaoYcpy470x9twMk96EaGhBg
zHYtDL4wSbGMib9DeB29+zbgh6CEIHZgvTAkn+sHNrA9I0A2xOOTfesch62+1dxIzVWAmc9jdiiC
TI7EY0ECs7VPBGvOj6nhLM7RJ4/jisGFQlcnY8azV5hLocRK5IRXUCD3NxAkjKucg8H8O/Ee8vPn
FJVNwjqcUDwj4cnYZp2u+fnB8Hiijpc/XlX+lqO/DPoYhjzlKaG1v4QkYQFo3Lqi3//STkZ1myuT
SEvfrmYX6t8CThzoWRyDdCEDq4UGgxj6QdOHPjZPTlsua0P/f065EPxdXZiJcgMZ6nRy4+oGs9hT
yOhwNWuU1s/hN35LRy61phaFq9YlG87E6hok9jeA8PgflRU+E3Y0qvb3KV7diadNsE4ODakllQzb
NfyEbESuovs+KB3GbQ4ZKV3XlI1w+wnysPfQfuC4AArXijNgm7z7yZxFOBl9+1gCMPOjXVuOZsFV
m5zWdC8mCNOKr8C4LgZwcLgHvdZxFDua24dEZxd+gXqS9ICgAXmJO1PjYta3UervgfkzFBgL1fAk
uV8PGpezaQGpkHTtIoikB4JgbPCbeUWYCQbPihT53xLzL/3cjsola1AoFvqQ5Q2bfeEaRXOnZlWP
HXK9gwQr0UdIaKgumCj0VroHOapC3h92PrtfPX5KCdImE8O3LRQVvRqZp1RBJpTvhSqujEr4QJXz
SDrQuuZlqoBqjLu5huO108Iv3y7c4KFFpCRwl8vewRzESiaZih6wnPgvujAVwz6MBpsnWJJU2Oa1
LVtejCVYJ7G0IamnVfEKFU3/q4WjJab48cGTEhOpT8Se+FDv/MDW79wvgRs+cqcWenKxkrfwRGyv
hBha3Xi64Y7ihTzETJHuR7laKU/hHR7vONJacxZLWgSDQB16EwY+YGCfKQkrJMRepslDQu6/7mod
jvVUytGABuPKT2gn6DEDRcp8m5vuWx0S/X7Q3nu6hZUcQx1Y/lImqCI64VwniydpYRwvgM5I4Ln6
c66Juf/TxMW7vnn03H2IxtLHWoKaKrhLshMw2jy27H1oDEHYAfjPMOUDQ6cC8hWE1OTOQwI9cdNY
EZzI656FJIEK5tSaVqgyoF+UB5h/Zrc/oRvpydTtRh8bLGWDSUKg4B6hgIVmR7oCV4OAK17X1lpi
aKMOvFO69Omadq5eY975MJFo/7ReVd0OeXzVQN6+kZ5qb/EF3CggiPiJigNvQVsZMU7vyED61N0C
F91Dim57oKnpRxCFtjNmckKWMRlw6YHgbw9dM/XaAzIbzak7F9d2Z70/Bp2Jg1sRE+5UzcXDwMOJ
YX/wMDhh8hcDXTEveOYim+z2A/YmFpCsjMgSn4Cz9pS2KPAlw3+kC6B3WzH/HT1YjdEmzUNFH97/
1nWkVCYzR+J8jju1W9dgoo8kggChdmbmm9dcSlGKm9JLM8lMhpc/1cFWwRz27dCOePm2dZRnfmfv
zzah1mcy7KZkh0nwds7ysAWMym7cHOtX2JOOkRG+YFGEpEScm/SyjHNxouXR/mTHNtj/ZWv9gqC4
s23FH5FYZaxJW8/uFQ5fzFGnlHQNdnLPIcEAE4heU1QfP2mj4glt7UmyT1UAgd+hbC0XEM3ZoerT
RpGrDX4/SocK3pRvE2Ce3nKst/UEkQ7jRLl5tPntBGPl87C4aD4k0fvgktxusUGdhAztr4xIsuKX
hB+yVB4HBXm6B1riz/EWzvXBFBYwb1pcHeDTqVfx8hAM1lPxv0OOByHbSwuho+k2GjyC3z+q8Tf2
dRhMnSSh3baZxBVEQLoSUJnidOOIeopRTGDdNa6iw+BF7cDCJRiYOZrtrDsCuGq/TXSrAhg+lPjj
7ubiFwIBmbnBClUeadEtVtm8TF5Bvsz/Zzbu/PK8KLsw98aYflwsEuAthDG2iShJ6skkQWCW9jSs
x+WdzzN4fn+Jb8/UX3ZDQURMvU5AVTNZmqEMYhUB+mP28jv/DUk3CdTFKl6TQfKjaDTSbSd7SST6
hOmMHnY0fYmQwx1ZVUdDcSm2komEdCWt6N+/uQ816YvBTbdtIW2QAFGVjlV7KpgVUJ0miSGw2lC3
f0MZ6tktGP16dNkJBFZxbKW5bHX/8AliLrv8YIBfvB2SufWLikuBfHl5tpEvkSRCjhv7pEbvoYJU
J0Gj/oyl2yOGs5624QcQQe9CoJmnIHZp7cKWdsyik5jSGJi3ERIdlofhia+UWOGLz3kyi65lZlA0
63m7bDD/k4a8YSGLfBABAOl9vX4LTUdFK5ZB6vQBCm7YnVpYamQinebKF4K/TnPe1KVTKFS+mcYr
TJHbEU44Xt7zhV+GDoT5ycgKQeZ3jHpaFOaJ0X0NwN+NvCHqFGyS3t/N/TV8YBL+YkphxGFnl/vU
ytKg2+4So9SG6Xv1xscGDpZINoGft1G0vJ92BFHMDLQw73rNxxuas+2QuNQrIeDVD4vDuEiLqqOp
g4J8CD7pgcRgp9vwvk6tOhh2uMVr/jGr1wP8rrXapRx77i3hFMTvSNzhKzeuf6XaheNqu0PAVwX7
W090b9DmYMQnifilPu2u6jmZ6IARdvFkT3BMNAknDY8z2JXqhL6jWbWu0Y8Q9pU0Qzb2shAIQAdb
WzGqgaVGrt8jlZC1GghM2IM5yT7rKvgixp4OHEU7S0FU+TbzS4N3Sgr01H84riCE2Bda0ohp7+Jy
kfW9KO+4AIkuoiwgiNeM3L/Gov+rH6/Jm3dgtiP/B0/RHh0RT5kwCK61fTIsc/Wo7taXS4n/hhJI
hdKoO4Go2oOSQqwbCSNT+TcD7j1D9GQX0OK/b35gEFvMmT5UALBi/egjm571J7gwxmXum+sEpHtO
q21SfdJFFVg4KWABf8hCVStnz4i6KdghY6ifIC7Rxlvx7tQfUh2ygWeDT5V0ckh+U6Jm4Zs2UC1L
wHwrSbKO5f/T7vWE6CGcQGB72KOSKox/PzKiKOrz5J61MFmIMhNeGqjCoRPfItSqc9aTUcVuym8R
3p4ymjDzKa0PR1Go9qywoAz34N3v6he36FdMR4mwl1mAR5alQmwyPvfh1q7k1SzdgE5enAMV/uJU
dkSYpueqpLJFiEqXopDBgFwz57W/wwsaL/xmqEs3aWxZXcmANPRoAI8OM9w8ebEKsnMf8CheZ9Yw
r87eTmadEDbi0g5Y1MwraRyNV3ulxErWNY4s4T63s28LdZegqPDV6AW2utCfhwY2TenwKlpcuIZP
elLbHXMybTjaRRFScdmxM+wGmT3MB5EvkWnm4AEfC0BNvceV/y3PbbNrs1202FVrhp2F+e47LDty
H0wXMKkPdt7xzxEG208Q8Lqr5vttu4INItTLj8i8K6OQg83f3VmxjbobIbtuWYqMhRGv/zNllOUe
svPVIhPuhNAm4yJJmf9smWmfwJq5YRrakXnNnlcujkWLrWV4ddqvq6ZTgcUVhdICu0QWTxCP88h+
CLcalNwKnNSAr9NgvDPQjC/H5NAigWm8naQE9dNxv6KgdKZ/KKaHjta5/HRoI6lJ3avejlWofcfv
eGZEOoDaV90N+chQwYWnizzgeXkSaJrlSjiFK4CoCHPyX3Z0of7TvLGhGT56/ZW05w2hXCk8KHyF
Iwn9Lt/OCAvWDr6VfFgygRWKrkZIBQYJFPSQWySsYY9ZLgYGeOjoHMsp3o0uzsfllxKy/iS2EXyJ
ZTOHvkBycGpQiYCvhnrbVl14Xm980AbjXC3hOOyW2zp4amoBRCWDKuJZGOHdtEGwwFEZU5D62lCX
C2qQG+tveJmIKEG/w8F0n+S7i+mgZQL4cF4BZvWjbcfLZ3sFOHIV5GvXm0HwM/Libm6jvOAXtvoB
XE2CBpu35OFEkq2r05quBuk4AIvPSrRnCz+CKEFk9UUaqQT9ZWmnYRbogJwDavIccCDCOzSWnydQ
adUE0dFLOn1T98bM9T6IvuC4+2JKm/DVr1Pgs6bi7+vIGsQUBhqNF5rpX17O6o3k2MBaFVdZRbpk
beKajAz6MAj1LCnL+p2ZIRh5Ncvhysd/Cq9XxNnvy9CY80Qa/wj6HV+IsGvpyTUUMu6wLqzWdl86
swUz/MZkWXZEd76/PUmiHKnEjl3J2kqJLWO2l/fU+5OqotVHw6NklaicpJ/FzUr3eib9C1pVIkUf
p7/KEHS8ucCfqP0o76skoMgU2Fv5zM6msAhl4uhVSI9BnR9KXQpJHswP5x2sNJFCK0JnUc2Wq0nX
DdqACVrSVo1wMHdG4yTRE2C3vntZBk6x7nUl7xKrDXpCla3v4XXlBCwgtvTwsBe4lek4pZsXwxid
Zm+cl3M69XHyzTuQYUBXy2ARTX+b2Vk7rRQpzzy1+88Mt3F61Mq5aKJKU+uWF8EWVYI/FkpNFYaT
ITT5rlvhquh92EdRV1F84pMnZP3hRfxk6Li36L+CxQayp3a8Vy2gjPUc2DjpyXWqwJzc0LiUqu0J
UCQETl9KJCnjvISRUvsCAlrYdZqhEBcsaZ+1QrNHD+iloY2yDg5Wfwbkgup0jpgwWZPSX+ETXm5E
CTpZdr+pd/XJJuCdBivMhKGL3SqCxkG3w5ppeFmf23vetiKpyjVZnMxTGrUBOeoX8NUrcrbEfurd
O9AN0sMzBlnG9E2GUEufkV3+yUdbC4+w+vtBO40hyNygL+JTiJ+mSSPipnvD2/nqhZWBJfzMi0+y
/OVsvLEmUJBXnLNB8EgSefYki5IPk6ZKFFs1MiS1hfw2nzLa7AjVvaw4njrfA6XY7tWuLnJoe8my
smTQRWqwVQwedJQ9lL2Fa6xeIQgzZVi8vVoTFHdpZtwo2YpW8f9TGC6xEghZqD5Xqm+0rHTJE2ex
QnbkfqXDGRYQWWuIX/VgVgDz4L31bEG/lWtLbDqJici/W8h0p+QLGhLzPoLCHbCWVtaFin2NqnSN
f95DVVtCm6GW7HJgfVMU9aiPnn6s09KdDnNv9TlY/9O+0m3lx0U3rXvBmyMSAv++HbgzuY+UZQ2d
LMiWmisA7vUVFSIb2C6jupYDKUKusBvnGZ4tv6LDq0/LWETzGN7d7VwljsYTa/+N9qFGRdLRY3h4
Ek+f6ITpI6jCG4SkzEo77joUpn6uCOOT1cL7pTKq9pi8xT5+cSxey9ZqmNC1162ymiFPpyO9c/3A
hbVo1jt3OCHb1U5vik03LtR8U8FaRIVrgN1srZqj/2va3W2yntWp7i2BHUVclqxyB6nSDJIeF77p
KTbrpU96jSCncbwNuqsCUPmLRT1kaQA2WomX+5L3woUIJjp1VCTGfXr+6YIELoDzn5w1iesGPGKX
EUl1ZDyTv66FO9vqxab9+AgTFscr1T4CRcH4HG3JWSTVLkKiHFvGiA0TQMNKjrRbpFtqPYAJ8Mdx
T+dI1Z8tpD8KqB3J11zdkpTecEz5eXymgLSQglh+myT06bo8l/Fobm3mJq5m77PntTJx+5/Qu0DG
AhV07ABlC97KELP7K7B7OnP+skSdZyD1WJuBRHMnBy9BgFt8Q9MkOgc8EenFz7wQmoB5ZsBOeyn5
zbcX+13T5bNOsTPYo/RNp2MZIM8Z3t6eUMRh2XIWDB5USqPa2dKnz3eefqv9iJGTuTMZg2TLuDKt
pfFsppj7wcrYaK5JyoVoAwcXMEN3ci3JKs1E1Vvipcq3NLXlO2jOjjGsh0S+T+G1zdRlUr44O3Pd
LZSBsUEirYxarUu+bhJhl5JH6EPKAccXtGPTMnWi5l04T94xcg6D3+pV3/qy0C2go3SpNCl8LPQv
dqYzBEqiFsicP0MfCcqub1/AIRclgxKILdQwRY8jquzBWGjaatzna8Waw3rFk+NWU/1k27IbKw1F
LdHuQVupEGuwlSizOm6u6L0rWFFs3GD4dfITnDzSlXttN3YpLy3A6v6wbCBe9antiKJRYzLykiNH
Tf880XN6hgmcdiasplOYIbgRBLjUJ1je6EacC/sEJvzDHFhY6ZWSQPVHTP5pUKkK+O05dnVnbWLj
Jjec+hjEBEaqlnIyqPj0z4GH8n4ABy+wv/TZFUHdMF1UIaaXKzN3PF6Llo3542ddssFCsBv/NuLF
cKAJU7eM6Kw2HZN+ELCng+MS1+20O5/hNAMPi6kHpRvSmfzh4/XJEOt2G4oxDlEi1lYZgjx0C/fb
vgdbKqX7PcxFSfJJyXc9uLYmpY6Icj0jlv/zpFzy2zoSgn9lGzgqyIJuUc/brOQZ8cWASjdB986N
+5V2BndAd/aRfL7hoRRcfyj3rRWNF3adhQgA4GqEtfJAFNyjJh2wM0YrlKPolfL7PJPK1GyHNIGy
AQiwxCuHuSj5JnW2p8VJV/hp061dHjybKL0CYhZ0PEDlMvoEHn9WCFx1asFk3fKKGAIy6jRDW6zb
yfWlx9+3GUZzrUuMPs0aIAlheD63ybEMAq87MO6OpI2UvUiyxK3cCKoZY2SJ1L9F1hoeMyTGWIWf
bOasfYvLtJ43DN5WKWh2+QSU1ZOpS1gSKibQYc9q/Ue/jrqXz1XwOp3hvHBHe0sHSQGCCz89rsXF
AbUJroLhjx65FJu1Hl3y3LAcoexeOrH4JTDLxqWKY950G5+1k7nu3etlCG5O7UKc+6Gba7LJvBv0
mTbj5NpvN2213vELQHEjxEiPiZNqumU0/gvo2u4k830C/stLBijJc5LhSaomUaSPbrZDalIXAL4S
feS5N7dRx3L37wV3YQH130AwytYQ0dekIi2YunW6towk98e6oMlCqg8pDjwVoL19ZmWgX1i01I6D
S1mUfqsiu/rwS1boaLEpQ3rOBkdoorbzWUypy0b/rJrI6VwBd+UcgJas2LquxOzd5pECPpHj/PsD
p/XemIK1zlSuA2WnX4FcmNiqIQLJY0GnRNDyhBHqa/mS9oZ4065PZlGAHvZW86YZ4h04rMMKs5B7
3O4kanhdtDg2MKZjcCnvqR0TyiiJeHcSYAU378F1vvGe5Dw2gfP+lElBehDBhb+6r2PAgOd+5MAX
pMVhkDq9gqh/Q7mOMRYJfazvn0HgouxcIX9XImTSHcFrAdnihhvbK1g+CC33ciwRUJqwm/bSxwJg
6iShs+dtzw/vH7LsVZLrtbeccUXjHHpPK/S7m5aA3cjg/f55Y6d8EUTnX6g6Q8tZ+i2u1cS/OJYr
92MmUdHjWJPj5FeBc7aTQjg6ARgCZe2RLgVKOwRIjb98Rvk/m0yjl16D2gl/uxLJ/KEBajsnKnG/
xWvyFi3IwhVZAssfQRuSl1VvQwdoEL4Ty4v1uDOuiqcBsleGwnq3k8ivwe46c9LGnfVtcRGD7yNH
rsxSLM0+5wWUHULUl8qoPSUUDHLi5by1VR2dCFwLGl1/uXZObs331/O3pPXadXSK1kcXNlAeI/Bn
6wNDyDug5dAI2Sp93eHqPh29HxHBj84GIWOGLcpwwHuNf0MXIXb2RJxjIJ512SvDlxbdxWdAqOks
gkt2Ym/9vSO1FXoI61YgAItcfTIguWQkRVSfi48JVwUBBAUjuccIojHe6KhbXaqm/1/Rpk3mz6Bq
Ih9tbJ2ni4FCZ3MiJyUiVK/xHF3P3N7SO+JpwW+jUCF6qXY7FotMOvw+Yr1acTco6D31LtRdsJlR
KhjqASVQJmX0RNYWP8GLlYzEh/0vPXDFcBH1eKVEdQ9AONTgoR1mwUGvhQaEVZ6oI+ZQg9HZU3d7
UcUFr/2eSuhbFXnGmrbh5e/iMg3KX/qaYxZQ04l23mXbcVQNmXBHSTW9jjqN7fwUgeVDKNzEsfJ4
gVz0X/+RtGsVNHEfqjGTxtlxm2p53hcGe+ipTBOtChDbEFuM3plA40J7xymlMBORr8DqSZ+dyRpi
tzLlSAtgcGLF0VRkHPrLy4DWknbLEqz/JLfa1r3t6Wxv66m9sde1lSwNodZgm9C1LUKNQ2fQ/vDP
XQtUQtq2QjowxmqTysnGsifm5JPcgxI/i9K8/nLCPmBRmyWoZCdEH3rNiKUdK/N90hipxI6RvY9j
pYgXGoTEUEXDTXLqQRRsZ5JyPwJ6Wl3dHzr3kPOvPZ4OHqKrQoUNpxfOFZH2XCHlIy/37HXkg6VX
IhQPeqZ1v9+MsHqFczBRzl+RQ4VntIygbWppt8i8ijz4r3aRc+K5ukWz63RH5CGpD8cRQPnTDsPx
JShbVJA+ZUs2Ms4A+BgprojG6KtFL6Ux+7/d1U5eoK2zQdNpws7J3lwCbuvjMnaB1vF6Jz8Nyzsc
gh8FWnu6X+k/7eQykd+Hsv/gyK9Q2nnvw6cto1FVEE93kW5K7lJrvRbP7/UdcwayeRuX78yWDOxS
Cyiql6f5NlXmlOr7HLAkSut13AJvzYkam+RqedMA/qdi7oPNwU/HS2yhCPrqA7GegOmSxrt3RvAu
8aeQA6nus8OpsL6dmHhTLQSd4qSOx5+rcssVefwVcjmQpimT0gJpVmQq4bc6wB13MmTi4BS87eSI
jrgA4gxtwsh4ms6CoDsOhRKsHbattBogDPYUBKJiygKLWmjL2fV3JTGRXdwcT7uiy+XKGjFQ9EZR
tzYkerM8/1o2DNBQzfga/s5lpZnWkH95ic+kkuFxXHi7v5GPZywJo6isFNLIlJyCzsgD7J1xVEUJ
Igpq2P6uFcHoHHeh91/NNTz0EWIPOoE9XZ7UeahTRX729OdAMFsv7NUQnrsziJ/CBUOIC5iC1WmQ
vA9k26rqF3bmYDSkNQankYe7PEX30v9F7W0kRFHUgvwvTrqK0CpabzZAxbgldZYxg71kx+EbDDH3
udtaf5BrA5Fi96+LLCVa2ZRTXatrEcVdT9sXpuHFgIrfxBTCgYe3hW8n0A0dR45Ygj3Yfv/vEgKs
VEGI50MbZgn27kBYDpXFpTynBmh/BseIqbRbQSPPUf6OafSlZb1k1hphoJOfZmMBIwFnRrqeSLm2
Crmd7TBKSKG3LF/1O8QyrszGTjRpVSUWAWMChKQBFWSFc84Abw3gXYDUYGz9mME1HTddL2ve3b/p
iRGFukmEWD6zdEu3Y4QWC/HCNO76Ug0fJbhT+yv2xIGM0QnABICBuGq77HAftDiKxGritADPQS1g
PukGSOVTNEOW2EDQBltLd0TtGcOAXrzgSr9N3OZ2RfAEijhtnq3BKGDce99AfX621LfJ+/FesAg5
M9Qo8MBc4y9jb4Sp0x3a+bcu0A2wPidRDInNfFzh6D95gX/5dNsWEn2Bbr26PsJPoBVWfEjpPW/B
uydGfDXcLRks4t23rPQb1iOXPgFc9PfE13o4k7JDjAoSYzBavhDU3g+yCuOcu7oTTGZrbwDFzPgq
qP0xz04ST1XcjZW8YSTL4v5gv2BC8cBzjlyaxjSyxGnwnxBEY7ZzOjVBm8KO6Pe8L5HzXBY+Re2e
wh/SHR4FUgTl5NqiaNio09Lv0s8nQZxa517nmMOj1uP1HZaWc2TkoOj7l35cxuFHIkda3Ij+trO6
kbYkcJC8bTaFSupuDpnpsl8lRe2Y2BS4juLYxFCbmTpKeS5Jd7p5Zn99ldkIlbXqkudg9TwPIICN
qaR5fcFKEXkxi4pFaKVhGEnLc3ADf5UQOEkVLH3wS7QBu8kOh4NHEYzoALI1LrccUH0ZQApIhEha
nZkfT1OojiUB+qi37d7cJ7Iyf2svyInkxW/GIl+u3rSFotQ4xizy/om0E0TIeKXHCHw41THaTcWf
jKv/JbRCUlKGYKsN1Qpj2xuecmVLAyqab220dxErus7AvTdHy2tv4Ft4mZvhuxWr/FiZRP+EBGwI
Ot/LMs9Xih7UxWcIfcwg5yoZLrukE7OO7NABe0/brkD9Ed5/kyj1A7BkNiXMMyoOT8VydrGd6xGn
UZE+hItce/mmzGuFVKIIdUFznzFFZr1VtrfVdqyrYUdmL1a4009vOdfuKhJjHbNYEpJMh1Z0FY0R
0cMBBHX4RlBsKFhxbgZg9wV2xs0Z3ltqR/v3v2oy+/9QGDXse2WHGIJMT56nCtjp1bLKx5maD3MK
Hc9wgjMSvq6emvd03Cv13Be74/Ls6WPetEvnIoTsiXV8igw0VCZRif67jPvmZ+MCqNDO7WCzRyXB
f2XdBeLEHDYoozcmAd2Os/ldoI2lgPK2CbNbgJgUtUryJd+ba56qSXhqBlWNXme28jvHm5BbWWtv
v8dqXCypMOhtJTubUCJKpuRo49TpXxdvca6X+527yp7hUnz0OutgpJRWUo4rtxBXPm9Kc7i8lj79
EXqgG+3InzJSQDFB++dcZpQjm+Hwy77h+tmrP6vcZXPRHegoD1DT1r7GgT+vJPHd8FJLEwp5sqVU
LFPKc5zUi7XW0piW5RihYINGyczQQf8olq89pbmnwiO5bHEUV9KpnzeUuK04l3xIUsRyE0GO9mZC
KDTd7XBcMINKdVfKOqIvTgBWuUBSe3hXB9qoJ5ToUcJltXp+8Kbqv1cOewdCJRFMkKgm0Dt1LfGx
vAimsSHVcYUavWFuNkgBr+JiR5H7meEkHa6cFLl6WN2O8O+B+tVJzqkW9A5Mfy0PTAL/vVRi8o26
FKqz5LxFw9dF1Apsijbrrs3l7tl3XbvFniYmvR4uNyJYqX6J4Rl6hYn3k6ELf0DNAHVfz3uN4zTs
r8eMl5JhU+hh/cHYOuILcm5rmVXXsBVf9U3iWlrnAqTs8sAyZj7PksKDO1JVZRAip7FSHpy+FO4c
+hqH7Lu2OSfbzNDi3ahNwehnKg8tF0gnJWALnhzfAWCr1/7ie9ze4B1b+sBRaCjzWCikA6EPclrK
BCBx6CDi7Uu6L8MkBpGWlkDOzJ7MQBf1HDpKQdcRZrDsYBe/u/WkgxR4NqMojFNouc3BbIgrdJVG
5wewprwYnjb8DCcf12Bnvz9TiGdGyYkVAfb5VauKTRYShax+bb1Rg8XtDHNC1Hco79BlpsDia2L/
M/3CC/ykOhZDCi79W1O1zio91MRuTIFfdecpfWQKN7hJcQvGk4hfaGy+/heKAWCqJmF1Zfjf+Beu
AUGQ2oYhWUbjDXEQOA3vAomHoSrkwwYu0L5g7NqUCYbGbREFZzWq6+Cd6GfAUgut1yKVkCxqsi4C
fgyAetjkZp6SVJMWmf5b+COUMW5hKJ6RefQKZpHaLtgKsbvkaSgJS8/qUTptCd+wLqQd6dihwhT8
NZGMeCmq/pqdoMymsGe6hy5kw4dXSnCVQ7zJn5K3aP9z3PgldeWP2XX4rwuQbOc3WD1dTNbJDVdv
A7Gu+sZIkVn+BIGXWVyod9A67h+8R4Bl1jft4Rv+u3+tknmcQ19N07xlzSuqY+9qesRTRuzuxkh6
Z4sUkB8xmQ4aPpJYjYVRi11r0KW3RsDi7V1rQZp3kRR36LPilo424m9yXCcxsDG8EaQMUzEXNKZI
1H5GMMTdg7HNvZcFbhlSInYmW6tjVxvNaP9hTw/Jzx4g1Aqey4a0oGqRyrMBfWhKN21tHDuxmz1M
ScILYn9TNbJGpqZ/3Btb0syM6qZDpebZ8cEy/dNCMl6Nt8KuZxPIqTreNs5/TYlDHIx/R5kNkRTZ
zNOH0E0S3BxYBscYvd19waLn/ofeYmJ/6SvRrRakJPL+BQ7PzbO1dN1x1lRbgpu0JuqyD+vvu/3A
IX7SOcRMbFrad3OvRje8+cj2N6pVWieo8BP3PH+u6tWinOd663pw2FQzseMAg17kHi/24rR4z5t7
vwXrb03ODliGa017AEXU1yzQ3J8qzg1avBczSVFCRYg+XoLNPX2FFrE4/kBrp85QjGqw0LQeSoY5
s0HrTEk6LlCwIZsUbp6gzxoUNkXE1XkRXk3C01Y7/pWTOFdlv+xz9N/49XHjumDoiVw7sf1QloRc
9STcaMzKLbSU2V2vLtpKiuttCWcYAEQjwndBKwQxEywWDj34tUvhvZ2V+novOADh0E5SmqC3MOtO
z6KCJTn9lyFmiy/cPq0oV929VDdnXwOxvWu9MXqY8gfgplDjXAaJITVoJnwTjm078U06nFqeLqI6
+1PJ3CsKjlCiSKP/LrL1F8I8/Pdqb+ZWH8NI7QQ9Z1lc1hxdpoQ1CwsxMqrHUtCwqUzK5fNt5O32
PMR13oK/QNfV8D3BDEYyRYCTSpfaODDKI75e8X19AbwfyhrnmfHc8t22iuCo08EcgQ4m6jUJG95h
HMoQgSAtQgt8T/MHRST5gS8LV2ooRfHyTc92Men8O1iY3UjOeNnOgDtSOrw7FuQ2vL/Qq5lTekIz
kEgDXcHpCNiQ1RzwU4z1UIHYFftrTa+1+cBUnEupYQbkMqRsiYWnAvEAedcby8/ZigrSZT1t4Jsu
LF8fa8VcXc5GsleTKOQlwA9nt2zgXk6cflVe5v62dN+VoRuFvrQ98y9Vo6oBDtYa8rWVwFW7ndKp
/MTBrA2ySpwxOAnlyu7SQXwIhw/sJdE25GXKf2D8DvDMalHzw9KfJGt1fIag/rAFMLCzFg2QVQkt
X4gK4G2cDbnxlSeIpsPABmokJeBpmSyX+Tffx+OUCycEU3YM9wUklD+9v3xMGaUaL9fs1+6VGnrz
VbQQ7a/kfCmxmpRRP210T0LxjoQgCOb4Ts7Hfq3RlTJUwSh6mQaOkXCqzcInw2EndWfZKyFFji+N
+8QacdC5wbl0nLkh/ov2s6NS1CxvMuKoDVEbVrWg5c7IA+ts2PXsm7TUV7LDIn/wmxFrA3y81kZU
Cmsd6VEqVnE6yv8AZPAaLbuohQ1+fyghTRqHHPCK5tnJgI+SE51PNMI9gmYfn2h8uWjYcAulmKH5
iA94/6N32gRc5BjdHeR+judN1Zl65uUjplw/UEr8wyWFEf8Lk4FJzqtVk/T/P0iYIWT+gqIcslKe
fzqxLU0V78HoUH8Ra+63GjMLFHvLSmWnSCeeu7O9V8c/AIUAkzkag8tu+nJGzu3ucCGAi2eAxGu2
50P+ThaLEG63t2gyicAwRW8lGr9gHe5zuUCEeTvnMX2OrXNMEtyQ7nzyFOvdo8PrH7+A1+ma43GH
1GscvS9uS4R+vstI9j69P/iScTULfhOnZkYOQFZHfMeefXATmAMhoSe82dzIpoflDsJdJ+JRgHRe
8XfCp8v4vSXgi9isA+CjHGUr+Eh1iLOtd5jhP9TyfF88g1Z55fcxy9RF0iwjWA5bAjihUGXn2rlQ
tdQ2XXjgdhdvZwQwSvi3eRf5heOdKSlB8ooddNU/uQqO6J/YCvozD1gTGdbZhuhN/DJXHeANm37r
J5FVd4bb93RhaUOBsKjnqIjVoVNr6aPcIpcw2kF/VVsGnUXCp7iDNOEcSk7hTvBA6OVq4YnKsve9
wfiEuDiAWwpo66MeVypjD1Oaom8LZrhHLZACUKyG62i2Rljg+rSKrtZgrrMANRs1XLDTzOLsfO5c
gbGWBaHb3VvjX3MdSGKwRQOZOZ9KSlGjSBnSh/t+NVPZlFWRO2Do5eji6LjByVHdG2cq+YSbDpwx
WxLi+S1m6CncbHT1YyysNpJOGHVWCto1gVO/pJFyJPP9XnlLDc0paPapTK6dacN8Aql0ab1iNe0F
GyYFp/k/rPPnjgOohEH3AtMoTQtem6W42PbVBpbQ9dsMLXvdSOt8k/Q3uezvqkmH08QzE/1f5xat
vWWcB1oScQwzJHrQS5GXCRv3ufuCgxWZ0gwTmF3Iu4LuSq3jtJC42+ZVhJmU9gjrzWM1MbAV/c10
gN6srl8GT9WuvWgrzVjQPrdhNxco7I9y9CMSJ58iQTdmn7Om5tSbclM/qO2lvHjzPcLZaDgFqwnP
fGLt25lQPixv1f5SZ4uM/Ftf90iftcR331FhIje22upe+FBu2sYbwsrTBwFaB/Pz3avV6McrGWpw
3tKQBrIxYuNzlAfOvzsGYE0JGL7hXa+SAwnPVYZFoeM6T7tB+CxoOEpSiWU0SE/tIocpjQsgjGsi
zejstwibtRY/LFqBdq8/y9GIq3Dg9JV7//+6WB9UM++hRTYxF6qRpSYbMschN/m/WfyT5cEbd9xy
VtWK0uSquGYG50dbjCpUaaSsPngEEYdX6jDW3ny+DiYGqGj0d2QUJH2D7kuNTwnT5N8beDcz0fYz
5f0Iae+NILhAjN7SeFmvklZyIVAIqE0i9eju5pJJ4xQn0/O/1pZVqyAGpdJyS4PvWHqJem2MsT+Z
bgp21TajoGxFMz+DTSPs5Fw2PFbHPaiSjJmjz0MLEVmE+JrjBiap6xOa7L9nS5Ysm/nxfrp2unMT
CcDqW3Gc7ybpkpcK3PF0p9RUQdYAK+e8a9oX4+2MyLBouKZv9tT4TNqFLd7htYgeliEzXw29B+4b
lgR/M5w5/JEkze7c7xNvTP49kOaZ4wGdb/6mWLtHEb5v5IiNHW7xP48bI/56mhFZzRbYcR1DxtTT
p5A+p8TAKN64gH10EEPi+uuUWJ0Jym9yofEfgZ0dvdo2NTsSnnnHXiDqhNyI66GJMniGdhEgqIsI
u2IeY8nKu0nUAKyGAct4yHnMm5jjYNV5wyUdve5r2SOt0TmVBD0HnWReeBu/UskkffP6Nju7f0mH
GFAZlnFOpAge82wYofk1GF/MmtHDMM6+Pjc9McS8vSg+m58NafCQZqUY2zjSkZYoUBOuT13qYIGq
zH6wGb94at0LRTIjXgF6pYk7MMLmHZPRI3KiZy7NCS2L+xeMW4NKvwiNbDo7+Ljkc4is7IyYbVeZ
a06y7EgrYqAG/6Rc0NEAhl0IzPJHGwfpkIGAf8saCy4imN4rUzG4bIadFhWbhh4VSomSqZbSlVqF
jQ+1D0IRtXC75ATQRGsGm0F9CYwmguUFxMS11fTCUCI6hrQO8w1nqWYEN2szB3AYpovGb0aRkgh3
0YRMU2k5XTLw5lB62CdpEQUwhToC7ZuGowtFZdGZ35e93bcZj7Wif6JC47DgmeSwlh/sahM1ehOC
9z7iroWsBApvRW+EtHiVMty0bCxw1eImGMeSoM5FJPfnh0FlZ2q903W9r9ucqsHh8Dv0BGoNC8CQ
msQEbEDdMccpaUihIxd7Prkft70tOZWxwdH8+DHpMO1bMakZiRYBDDVcLRp5twlfO/VIRf952oAx
QF64z0bNuqajWMBLC4hMxhYoXcGMwOmSXssaAvPeNAcL9dtkcGVBdaipuagy4oUpQFe2X8zhEJkI
VDXPbhAV3ALqtjuxYP3EyMVeyrOR31sEAPCzNIzPMk9aE4P2d/R+TSSy0H6PkY1sJodg6CZ0ngra
IyYxUwxC+8B3vHLa6LkCXzKmpkMpXqVDXz4WEv9OuFApm/7NCxzytVWNkNJOG+KgXB0079dDUE2w
PlQYvlluJ5xPLOVrXMn2PefYBQ5rX5ZBHfCGkN1kpQSFOcEPPi9Bii/4VN6IibeaODJXsTklXE4p
a6q7FmxUxOHdBFJEf/6jSH35Z7HBaCzdz7HuQYzwQvY9pJu0xnMxbAAu4PvgG5Ifs1h+ndF5ozVf
fgzI2RGu0nsEHvOfvZTYEjPfMKNJRje9bIfJRDvbkGJ1ZgufAdo7pm4PbuJE2xvb4ubuSrVW9oqH
xKnRB4TeVJNA9RZ9vsUYx/17BHrR5qCu1s5hj9sllf1Wg+xJAFENKmqkOvFoUGIq+y9mMaQUI3Jh
Vp1KH4hl7MVb3c+B95M6P1xKhEUJwDIMx9BT/5LOQt9wMU14sHURWT43abWoYXH7XWtHGTFCVqpq
CE2yQKGgoUOTWYAiiQZg15/LEfcIiMAl+aIb6D5e7eZwVO7/bCneFthpv5C2ke8uvfoJBDFS/98W
i6O9CiTbW3pV1d9+CjXgOd+oPw8yn3/eInqkGd9KkOipseLOVoDdVFI4OksRxUESJyEpsC9m2D8f
S+0fN1hpucBahpAkLhtnTVY74U8ZbowBnbYK8+R/3Pl+LOXI7rx+EUo69Jup+TIxpimwAVwn9ajt
m14gCCD/un1f7ebZdiD/1NryxsWqZA2nMSl1RTSm+rqnTsmaGpMqD/giPZPJOVRPqBQhTu38g9nQ
xa4mSh8bqVEkyGcEHQCDWknrl66PDEKVRUoyhuzQ+Kkv/YUDurOulwYa2tLpnKV82cPKnv8Tdb3z
F+gBdy5gXfAbwwc2WOkw4LRjGRJqUyZ4w0PANFdyRbDthD11sFdCM/OqRnJVhhtPfs/uA8qPyB3Q
hdh6dV5A1I4JUKm6nmEw8jas/5hBv6vMs1zMU1np+4vmAc+qq/wh4+4Yt6yiympmcl3HfheBTwEf
wuXjElcOmGZ3UaZvzJU8jN9R44x4WESlymIO6mXuSn10/Uo1f9ryS8WhXE9RRUDX3yoVPyYumwA/
w9/oCT0/FWvZ2ZpMSKALNizbo39pSSEnwXwGcle97tlrKiZfNZEzzCMDGGW338MLJo38bs/q9ae/
hKfQqc3HSboM4A0xq/j+rjFeYZ32OQ6qRGdMxIVOa/HOL/kM/AhmaENvJ77gJPNvR0wN2dQ3UW7w
RD95IIK1C2sKwEG1CbD7EZ8Gz8S4UQH/0WoBOBpaxvb7Kg1Pt6IU6y6MlVnvLPghuXPN65ATFRIM
Q0A0o8D4lcX23IW6B+UGHBrnfJN9yZqvlZKD+Dvc5OB2BumFKQhFvnuEcq2MUIL+2ZHEQHa+PoQf
xAJu7w9RK5if+BrgkaMT9GTaOMQHx6U/Xa4aHqjHLw2epvYlQLAZvbANWG3Px/WWWWFk4XX+1oR1
dOahnCCjDXSTKZ1wyp8zqqdH3M265LjcX1QtZ/ga9BO0enCpS68Zr10GT+ALGfccB2m1OBjqniD5
wYniwPN1j4p3CkPOawcTluW3HWLVncfpTtSer6REGH2ONuewLMzZx1VS0Xr+0ewx/GUaUn1D78wE
dc+W1zZmGm0LHNuzaB6kOKrP0j/vlr+HkZ4yOWLXiHgUEyRZMjo4rLnd1tEZtq1eRvtM5gaDvzUT
6J0xt6V7l+DuAJBGWY8ubJ5sIVj+pVIy/uXfq8n3D3Y9IxWsehMJ3yTa6rVWUQR2qXkv41nSN65S
qsmzWrEDdoAVm/6sKWrqbBI+JcJY8uMHnDafUNCi0XO7raehApfI2UePBw1tTjqzC4wkt5cgzcGm
NlF12Q8oSPhugr/okuc2ZwS27+drw7XdA2pg4g8ThXpsWgg8LvLWeODb6Xr1D/FdwYoasWyzsg+x
C7Y/QX07WqVMVuZTYdNa3/XFeqtpLGUUh7aFaD9fdUTjDK2EPFC3gsz1CzxoZzW0/Roy9XW99Cx2
iLsCa2+OQOKrbxlgyZ0oIwK+5S3cIxZt+vuRg0UQ2spUBxIkEeXdu9Kn5s+y2yGk1/OmTgO44B8w
sukNlFN0GU0h2ld2WPflJsW+C+YP8cVYnAkIOmOOR7oRlWZKbPaZxk5aK0Im/Mkl8j6xZxzdplcm
BlN27DRwSpkLwyIYAWJk0CidVpk6/2XsnTVL1PnWxVB3Ybl8hHbigHGsAgJeEm1ytb10xJzoFgh9
vaMO7N9RBDapeAlju1yCmAQTCjdrcBnzRqH6P3mgYXi33gpyT1VoLhvHmfzTvV+3LLzyLl9eDYqZ
e+l4u9a+SM4npLE2OqKRdf4LMmKHLOYA1nNFJWrQpmhaCkYmJ+unoBr6C7Q3KHHPsdnAdRnTmSaI
rtH4gRQXHesBRbM/4kiozn2ov0zN9fb0PUOp6a/fwHfjiArLTy+KT1HqPu+PkcizW3mCmqL0XZne
VZCk6lCqVxOKi8/Xr1s2ekH/EnTkAKwulpJE3TWcUsf9jpKOHaPLKkiw7OsxXpCOgVeGr/VakItp
DBO+M1U9LSBxSq7vBOwTNj9tlukRLdf/ayt6h/q+ORXWtC6N3xB4vnI06aMrXvESasQ83YTAdCxK
CGfbzM7P7en622bu050j9gyLEmCZdbEHYksrCZNG1hqnn5x+xN/kcq7Rn3jtsAcl91Mr5jp7C/d2
ifwILyVk0ZG5i2YLSjgu+1zqYhT62N7NVNfMFE3DdqXhvdXP88Wh1ndPnF4Po8QsLd+sLwRXVRkn
Dz30SIwG5vTbPq70qDOp6zQAHKl5OPDPBbN+6ETAArsII19Eq8vBTLkVsVZXmWkZYU+8bd3QW4it
QE6imDFhcpwOK/1GrgFxY0cnIBKaxc7TZ6MjkoKlwVDkKuPHnQS+GgopCM+kBwk5EoFP0QQhV2IX
xOh0iZq2at5LMgFh3NQzq4lO/EoVI4pqTwSD6ufTTqMGybbhvWylER30P7xxWOrzOKc0MKFPOZLb
0SAc7boPO8T5kle/uI9R+0hOJBcvHHF9VN6saG/JH1Qe4F35zNnPgxK/FMsN6SOGHvvGUUG7R+wr
l+/QAxDWQEQN+bfzBoB2geujXmzzBY/vlo4wUdFQZ4O/RfpjcbjSoNNVRRCfb+uhwQIvKPz82FZA
61YBXX0Q5UtMOcpow+lpkvxjsmSiirD0oHswH4RxLYR0gkRnuAuFIlpEaQv83hh0A8Yp1ehHcAFJ
zOx/l77PogkHKQq/bvvurYvkmAYFE6HbYOVo5HESjVi+spEVNjFHdR170lI1lyly/WCd5XeHthgx
gOuJxvQuhB9IFj2Hj0ZOAlTQqxVvqGGFolyvNcjnKHXzWJjej+d30vVBWEp3FYtYLx2YrJyqDFyv
RNOFPCMrwNhyISyvegPA4c7nR7ffcpWbKwp0CMd1SYAR2Ww50pJZo5OBFY6mU0ySOc1tlgbMIOEw
+jk8r7pcqV21BXISMCfR2CHHoLfU45/hONxHOxz+Gs/e8BQFLIuGOy6LWc9oFjksmzlRAU18Fr0v
eDiiiJOIphBv+kYd9sjTR/Wxxa0+MCvV3brY8k3Bu8NW7hf7qP4ybOaVoGATTf0WnaOAwtyn6fhL
95H45hUPRfgGbS5YHF+3SPinxQI6xMRuaep0zmYI8WJo/bhdno+h4h2g2ObcF+E1LE1I4EhELTWX
W1v3SfWMz0+DJVW5DfpVySHOdtf7IKenq7/OuhfH/hj0MwyQFEyNZrYkmNTkMlE2aoOZkV8ddA5M
kGwyZYstnJhMOCGZ8TX9KAJI7YUWHQgtlU3QJOMn9BUM0PnZ/NyFTpEPoZidwRnTeVHy0/DL5YZt
2wl/NnNzCiHWroE/kldUHOw+a0ZQETXgfwU1i/Sj3WXfipmW7sQYhmR+wHHjZ4WogqbcvxHxF34b
5Jy7Zj4Bi7cwzZ1kvRLVJ+XtmLCwc/0S+1pORS1dlNM/ECJLpMUE1YZz0z4S9xHWNGSSNTg0NSeR
f3CkITqbWseapE/6Bzg/W5l69eRaZ5ow7G/g4Fd4CkxElC4Zy+qivGJcCsKIGAY9OqcwwYNuKb66
GtGIMyZAoB6gqFE+3vuhjvGO1buMBTAAGz2H/724fwsi1NArz9KQ5SY7PCokZiosXxiveu3BlZLH
ErEY37FPhF55ceNM/cO9wMDoTRvnxocT0GsyWyqdCF7FHQzSv2hhXoa/BUv7Efnj1pTPhGQ0/4g/
JVThTPaDo6AEsOOXexlQA3A9pO1l5smC/+phkxZKWvAu+n38nGlJw6F2z+Z5UUiDQWNEq5daMnZy
zEpHHM37q2qyQS+jjSjNY42PAYTTEfsBMu/idO2Ix9oWCffe779MQOvC2t9AFz+kb65aAogZ1SOR
N6zm/lgFEK92W24fL756JLPfzUDWRPL5lbKAvlfWKHiVPFIXeRlDAkCcK4FL/lTHYOMiVmJzJ5ma
/BRMjIP4EfvnQCWZS1c1c+r1RhL0Ky5mAhihhdO0vic6AdZUmYAsTgqTCvzpJ2naKl5LCAaxQTFW
AVkEJYNFSW+BTZyWcdRhI4icB9OW/m30trYZI3/LzEIMzQEglMCwpFQUaZZW1mY6d+8w9/qZXzfg
o+CX/dE/cwyiGh+qTXXdZ9YQugcdxLJ+sOd5/A4W3XdEwv4DUiuyjgska5TjvNnTh53YRQTp4BZ5
7rpEJWRgxWPZBuYD2K5EIlbXzo5uwvxHh9/sk9o9kpW04ENUTc7mSOjEKZ//kXPEwnx/uKVBCJhM
pPYRLafQY6PinMFJ9tOJnQVhJpxHJR5GEjkMbuu4gRshRRtlHhH2IY+54RpVCDvqLm1bPSXckFDQ
v8N89WCJFVN17az1vcnb1uEKjf7VvPfwQV7ekXCuxkv7waLpJ75wmQOGUXGWHsXAyfr5ESVSi/C9
SpFkfpjTRW5vsnAgNIUcNmtuuytoozlcyaLHpuKs8LiulZkZCzIzk/sCTolLk/rM6LeVUH3clC3N
omr3m9nlM2Ay+pyod7C+6HX83RY330t1BecnNPoY4pAXA4PquaPD1XiJj1WLoqcqstrg21EqMlWn
4aUugtWegSEb17nXncRCYjF241yNkS6gUQq9pkAwAmUAkvpEroRoW11s5DxZMUnCiIb9O0UJ0JGs
SFCBnHVPVthUwx8GAdn4ZKTLAIrSoPVK2QTU8+g9iqZmL1ZFv05k3/PajeA/++B+ea48+rZ4O+qc
JMZAUDiaOnRur0FkzCzioEltkD0H5Vj1m+cGvIXYsAeXh6YB72X3QykxGOXaJFlllyRvFn5e5AQT
hHAvl/x0sF2tp5Y6NRSkB6Qzvs4/wpUF21wlr+masf/6OmgQpDDnyLQvd/xCkMwytfEGNrDyReO7
VsOSk7s9UzFXcIRrytfRNEZX2h6e8L8eeckeeSaSqhlnUxd7W1tD8vPAIMQWtxjX88Q2eEITtz/I
bsJbE/OL3T3Jv9mOiEBUTh9op863hsGcL76GyjCXTw9T8AXUJqhjWhtuFp4GN7IA+DDrgrsqrR1k
yL7+laoFoq21lzFnKy05veGlBHMRAI1sdeM6Ikfrdhw2FqXmst1CKKP39rYi/3H9NhVYR+vjF1Rf
pxlgS/DGV8Zlcn27xve7xfUr6hh+YX3iXG0H1J24tPRizDNSf5sLzH2TygI4wnQNQTvK/9YjqUNf
wo+O8YcB3/rmi4+ETjXNlU8oelRlRQkJA9pMVDoRWhuLS0se83jrZgZWqKQu+XdbBkG4Jsfsg1RR
MbIQ/36NFX2pt7JoggdMjL2V2VDDT/VcC5l6dAglSNBsinywxqOuTZR4FCzXWT3/xVUc2v77DEt6
ftIx+CHrYP8fnpiRbwEvm2D7Y/VVnUa0AsJgxuvbwgbqAL46Q4wL/nZTboBe4I83gqByh5F/jlj9
xr/LtYiGTQvhXzq1ABpPHbjbsi5bNfRrBgoTThxBkyL8oNzQBvUAfgX/eutKMqPafLtpuCH5+BZA
NO47OhL3vWUe8pqcDbRlulhUKImBh0Qcj0gxla9EucH/7N/6Ea5vzQECHQ/79QikSdpDSImhFr/M
YamNfoeNnpBXLdYJ5p343jCEgrvSWv8ESOSmrji3VceLcSLyxrmpjn6okmXylsGA+b8ZcZBSLQAt
olkPKrxif1kA1kAds9IMaz0ejqbBnGFs+kWyYXuuyKcFaIKhDxLdLjcznEDkM2xhYE+l1ugKdpzO
V9rMwK1GBl10muFM8JeOlJixkajP0tVbOQUNe/eUiXNXACfIWVXV+2vJuoBYz8hEof8IIZ7JsDUT
KA/QD1DWBUwAvVpciUWzHo6Q4iRjb+mBfeN5KxgNbsVD0xdjnzn16JUUl2VuPQuSZkOV0cWLAavd
AczKC9h21mHH1TD4HrfuAbvBlTQ3M5dnLDi9Fv/MM/FdNkoJfoIVS7FgtljeWOD0pZgOsL8XB4UH
znnAVhSVNOwD5+CGKXXLutMbIQWd2ERgAmHCZWLxXx91//BZ1ipyGG6Wb5ykRi3oreoelJ2HDKVK
txaYigFFRZG251BPF0b8tDNH78Cmi6lw1beQ7xR8sILzi8xCZfJ1rTLJ5tBWqJNkCjAOQCq+n1lJ
LRg+PO1TAh/gy3u6BiCck6SemkhJq58dsPgzBKp6GasqcTmjEjnZIiNwLMmxGwMS55UCS3Pqc8qU
HKMKoT/TIEwk9iauNDnRVI49E7WG6qy4H/Sg4yd8E+PUj/j4B6i7BDDUGYpDdD1lUbcP/SB3rcYU
yxVpSZP2bBjUKBu9yMtnrFExp5TpPnFpl79qvwGX70wwuX2qembsvKkOP+2u8t+yXoP+/dOqMcuI
q/7FTpDnqQIqzDT2LUhhkkRYmWDVkkrkHiGj0knWSxEw/WcLwDDJTjToi6YXvOS6Ah2sT+a9sLd0
sgCtSCaYzgvTKZ2aWYnXhzrBjVwQnZPYXpYIdd8m4D5qU87j7IQonONwWvTnlHPLzxRt948/hq4H
9PpGUCgDpULo4Qd6jp3IhvmNckRH8GgddRFXLuXzhtlskLgLHX3wQl7J1XTHIUtNBtejeAoxIT2R
QO1JB8GPK2aBBgchYdBTPZDxDADTvOEEBxx19dge8HRGCSHR2KHu/DqXEIWvLC88nNbHAJFs3X2I
8ecTckEndTlGSOAIsQDtQvhpZEtv4kG2OO5uxHz0XVXKdf7sBzwUmiX1Qy98mXK+xIseMEMfuODa
EwOFv8WqaENJNNqwqqLQ2YUASvh9vWdpfHCFx+OiqJgbI4BAqdeTSU2TNnFBzQps7LBQrAIXQDu+
Gw7Sgb0TSadtoxqNgQknnzQ48hLRj/aQOZw/d9nxg4ieEOuRvcYvFiiqXPsbz4vGbL20GQ5ZMb95
Ya5osRFxGfYbdxnvIL3aZ3oTEL6Li3RLda61+EJwuM8xyn9uMLJN8sR1eNEHzcDKgx6usWuc3iAg
JJQTWg+0Bu5ilr7P4afs2IgejUV1NwxpV+3cjr5vAEQVV1i6ZvDqypY+2R39f7s2EyAgacuSBvTE
aZNSeMP6rYZSI6rWuCGhWqyrDuF9zzpn7Opq+FG2oDNZ4MWS3SWA/BtY0++4ZRw1fnUWQyqDy4pG
KXgKF4Rsz23cyCUsHU4X2JzajjznoEcoYVHflYYi/ljHqzrXxTAJHaVNVF2iGxQ4ggpwIIbHtCnv
lAVesaIzknlytZlkH6k0ZNKtf6G9DTqjGq7Ftl9BRh8wfZ0uFtz+4htry8187EBQnRX8GFi1jitZ
73zXXIgv+7iFCBZtiK4GS51NGj0jAzYjBwaRh/5HlxdPOxODD+xtt4/7hm+b4lpHziMcbyljlZIT
oOMZBygF4Gx2gJtnBNogOJRveOp8wHnNYjWuH63p4EDFTF86O+FVLxQRoYI3w2ZlfndxOGvWK7kp
wTGkl6IXvhMXMZ5YPDcsXryRty3EydcMduD6ueyAvrHA1hABbDaBxGd21yE2hWm2Boeyi0EnK+fy
f1owIcc5WeZXOcBHmaoOSclxIRvsJME3KI/U73WwzKW7WCAGRY6Bvag+D5nL9m/Q1vJsADSu38zx
NdpThQetJIMzbNb47MSdiWXj7WoLxk64fqRAmZMdG4FQJH+VPxx5FcgNGSfgOxMKF908abmBLRLx
UubFu20m+fAONshClNq15OgdBScMmVUnY6Yb/am9h2YJdWy4GC6fcHXPNfvVeevRum+ns/N6SvDh
diakQ4u5IiN4LCiqq+lWia/87lEe2CUzl5PsMFDE5XeIuxxHwpSmdzubZ4kWRXzE6NQW+HTWQk5u
SFmusT4kqYkU+3PGjPThPEKvIt1CbX1GPj77C1O0f1q7LZxlpvH353dqgUH1d8lsOR4rSzEfTzRC
vMRT0wunznonNw+LO7H/IWLPCos0RmYYo62RT2ricIYv4FRpO4skJ93PJ3idit9Sa8WNCs6t3CUd
RmrPokIkRSYN512Xe6ZExAp5f2Y/oXa1ITJZpqKAPoIRR0dTELbEPcjAzwt5YIUZwl62oFdwSjso
wWNLVIjZsx6lwIAaJ4q/VEG3QhqdL5x4lh08hTHVY0wILRBYGNVxo1eGV8+nnwFb93Bs21yRBXsW
9yQMoQ26WJDipck0/w/kmNbWfKC2L+Aw+n461VgVl2oxj+zpTfEQddUZj8FE6bjsQFeJd6XVwSd8
jvQchlIogrpZIP/+jQBv4FgJvq+0gBjGUCnGOAgD6EDRTYb6DeiqfespPVKTCRHjk+frwkNhhgcQ
xQmSjPX2mdjHy4Kq1LdKDhiOY9+ghd/WJCSud+uHFedguvBcSyaJWzpI1EJIfwD7SKY1djxldYbu
HPcEzJVr+BStdu1zjs42b73pe6SlYJ3S0X5Lj+G59p2qPEgH/cOZSMcsCzeCTzdYIQgUUI2OFhl9
x+YfBuZEsIc2jh/b13f5Jd6wrP/E7qEqWkClVknuJLEgaDKm/vsmXSzMeOEEU1Jj940s+wkO0SJM
NjZjY1TrANI1NCiiF3zk1tsJdurU//HBzPd1MoGPeEWDUfTe67av1K/rghqjzHg6d84Vu0IlL72a
0DyOWRJGqLs5VpmBM4iuB22QXMd8I1zWUqhDhlijpTgoj01vb9yfhGXKZ/8HELOK2miL+Ftwcd3L
O0K4gberbX7Zqzw4Wh0iE4MUsV7UqR5IYuhAfx1jEE2ISRXAayfhrjx+knUYQHK6Poxjvlj9GrSa
FlPcEoNgsKHOd52VKnKLXrQ+dVxjdo4TCUl/gfbjdnYu2Kg3/tqfb1ZubJmgQnCJugy4oFtlwhsB
SwHDNPMwN2dQJdGXbFD3BfsgaPrO7I8Dkc21GJGLWlSKzmexjHPmkan8vot0aEGmgxwe55o7hpu2
xN3lgOQbSw6EHk+bVxfYkYr7KnW4zLFgZbAo60kFc8NS4IwpTMMw+pSazGyi8VIQPFKvKQdlLrDP
pnRvKWRDFfy8IKxl3BbMwQG9yUZcc3Ct5SwsJo8HkhufAmdp8tuGZfsMT0bieIBMFdpVZ8xFuE52
Sr0HCNsESZt5vwIXTMgzRdcP8Wa1b2CqL5hTjpIo22D8iG9z59nHRx4msy0nnYLL81FBwQ+Yl3pT
m3JdpdaanfyB0xx8eNe5Ei4QcayXi1wl3VVlTX6edgWQMMFkEeDrAIbWWQUHsN1Yu6JgGEPTh/oI
ww0cC5JGbnyDugKGj4Vqj9DxoLv/2vbg6mmes09dv69TvceUdwIUXaWMyewsv12xB9XvingWQS7W
8N+imcH8wASDq2A+MDkXiR7rUOqc0A5s48ZGR2ktKfQSRQiNdt4SMr/q2W68IjL82tOZ/mf1anoZ
v88e/Wx6+NPuBRltr9KanxejJzHrJfODugkbvQrEeC9x3Xtzmq0Qks6nEBCV9l+uizNSsqSyQmxR
vD3CN3m6bNnDa4Mn4lsnLrMG9ulVfewUylUs8wEo8k7QQnaUgZbLVNXaX33n/EY+YUYxcopoCzYi
p4XNEND2VLeZfufCaGiGzvqS8W5bRHQqEC6IonxolH9+5+L+rnTRwmNuUsuAuI3WNz+97JbukGUi
EEd6ymNaByYOpb+7FR9cRsPs+DKOzL2AUjWg3Z/IvhN0q8pQZkJy/j5Hjh1ofPYuyLl7yhJ9qb/7
2OvbzjXwdivw6meY77KMA6vUuc2aZRtkbjqNiQCm4ymPDyWfRYip8YqnFN2TI//9yqdCSzGtZmqN
A9sCvFFVI9jSRFqEeC1VfxGgh9NNpKRVZ96bpBOc6l/VgE58S8z6bMW8QFD+1gxUkhy1Stnc7Ry2
/576qXRHXuYfGbfZZ+RkCqtgkD/3dDq5lQ1V/Wb4qA7tmnQQ1s1+zU+yVgRse0wG4118gZwa9j5t
3c+0A4P8grVft8DO/OZ3YVDmV0uG1GNhOva1dcRS4Dkg5VSsXgMpgJNiK4LCZerAWS+vkgSDkq7O
01bKexVoQhwID/YowNShnCTHSEDo3dQ1WCk2Izvj/1UY+1ciVgzr/r1wtK8P9lFvEFIuWiymsoO2
2zZ3K6eAJHMnu5xGvJWymQxj6iyEoBIhlnMWXqqHoFGFKtB8KI9MPH2SjyGLEjW5mm56AbR7gL/L
hXbs92bKNBKgH7Q3RarWry8ngBwT8I5tf/CFXtJCiUfxHJOD7kn4tHv2iDdEADULhRO/Mo2RwXzf
+Iv8favupo15I6EWvpJ6vAthgkkdaAqpbI2V/Ug19NbsKGVBEhJoCA1w6yl+7Bhn+/HbEugLNHwf
PJO8dgoUMKRmPVAoeWUCeIdduAZ7t8kYggOAV5DWhcfOexgvLJ/hMErTs+Gg23HBLCkVPbRoLmw7
xjbLW0uliogc7EUVQtBKNFsfnj2ka7JHRAjJNiJBTktdVQfgVAxXvXLhDzocu1a9XUi3JueAqPOP
d/KSm1qUEh8sWEtjNanTKLcSMSto+BXb21sTLJgyT76iPC2zZN8FI5DTSKNoreBSox8X6bJEFj96
fIBJ0gkiqBBGXhVatOWdXzGnAJBDg7efNlMBGUxumo6hMA7lus8XSHTZ1wqUY6nSg8eOEVcmVrHI
3DPk9lpMZZaNrs9M0xpQtlRrHVMFmzOlI3beiJ6BV5PbS7604H+o6o8AVeksD08Xh0kBWkp4Qf0q
W8mYhYFC+c6ytGp4PHqSrRr1C4TXqmGIaw+1n7JaSfOrFPn2176d0CRavUBcsWcCzeNRwknM70Bc
mEhMxCxID+Qzkk9kMCksTbv5r0IA8Z4nIVby/RZ8KRWOKfLx4bkZjd6H5BFsoZ5LEp61DpDc02hc
3IRQRcNVZUPZVpJMlmXSJRONDJN5Zq+soTYbsBe8bMgyu0xYxgNPdDSPB/ZkvTZY3wqv0oKEUvJa
TZa1Wp8NZ6Z3t4P+piTSWyJxKb0QeSU+KMtQX/7dmY+lnvhllGto82XMW8kXnW0RjCa9RtYqTiWl
KjIrd4bqD2sNe35XlzyjEbDtuxkA1i2HVd8gk2ESjzE6ZmOIiip+Cv7YMdp2hEJx9KaN+cjkrG1x
Zn6SMfA3RZPDr1ZXpRyQVUnUDjr2mSpYvRuZoyZEMYuvv2HeuxaUtB8rr7f55hwC/W/POgcnuZ9/
W+gdZCNIc2Y4hO2M8zHa4FqxP5CHv9H8a1+3qdIwrXa5jOgOPof9DXiLgMMVAcP/jnN5OJQ2JS7G
0R5laF9lImoWa04PoCoqqk0Sd6sd+Hpo7M9mYxAME4jWoJzTpzCVSZNSbU9UZjfdLXsNmecJSDi1
Mjz+meMe5ltcbDaNPu8kCABMGNYWd3VNX3+at/G72w9NelATbDZQT/13HQ7kizc+dkEbLebFvo3+
NOUIAi7GumrQG5Bo18zART/alPu1VILj3xLAMLUzUI6PviE6T8wlbPHLfxrEIO+k1W+ntECkO2WK
azsoPJ5W4F4zv9oS1zZR8IKtSYfWaoBueU3bYJAV9wd3mgu5NDRKM1cdDF4/gpWryN5CTbCXVtA3
dnYUQm7dmewvTwly/lLE7xvNzqf3trx9nVFpGQNCF9vwExp7XC8Ca0qovH19gcdX1kZ2T6zxuOtq
wLEkChss402IlPVy+2kYWnBii4Oov2bKtwkGQhHmLQ+QeK/11UE5CRkmbxY4JZUUiPDhM4hHhtrw
IJymSYP5PC/BIVzEq+XkANZnrgNOdwRG7udA7YX7cs4NUFjl9MZnJeL798mREDSZ5VVxe1PcrmAd
DqUZhJyma06kMyRhA+EJmDiAdhCKP3FMojKb4IV24Qtd5JaN5kL4yyV5cnnT20fIn63xGbMDVN+a
gnfzFLvE/xNavLSp5xn4r/6bPYQBL7ooydwqEXVVckM85tbc6Bflsuac2nsNVaf3Ifp90EDwJkPw
inziVnG3mVlM31ERV+N/g9//DBn4gQVLQx9T+WQkGMdlYlbuGe0hJDc1shC97QwfFeMcaEqRUZJJ
6qvA59lhKZg2R+200gnp1bcB78lWs/gXR6WvNdrzAph7cvlXYH5nDzEws/SnVRxOjoduuIASmg3r
t00BmnwyWOM8ORh2FF4D+7v2VAiUOmmVvfCH0oH24wmg/MnOLyH6Ne2rTkdF8cBay6tQZXZJfXuX
+Sz3Mn4Dh4YFxHt8GJAZQAvPpO7TTCR5R4iMcqePVulNakWnSrFlZwYnGU4BKQkd6bN+HgIPqwMM
orJqg0BpQAoJExXFk/5Wq5pDwReYtzH+mYYcYUfe0Av/PdZ3FQ76epgOYoHi6kO/mnJ/g8j/tTdT
rZuxLxfYepUdht62WL/ptWYR3MBQUfhbpwsYhIQQs9UUR7IIqRgDuo8ZpxfhBZ/v7xdrghWdXkx1
iJQLp6SRocXvEQGxcJJPe9kLi7ARgRYg2rxJMRW6/EDGXM499u/1+KU8hvGcOvq+nb8kU59qbMIL
G1GrVFxglWBw3hA35guVPyxRppuOe2qDT1SbHVz0/UZHc3CFx2qy4SQSNp5/4Er+tWZXTzjybQ7h
S7QYfwDpDknZolssUgMh86g8ANBc8O/G7IuTOFxUFT+oR2cvhSsJMs37hVpUCZubOTLi4MhIjGwF
A4orj44HTZSNGwA1OEYrsPCAe/tmKgxM07YLMzwOtT3vg08KC8/C34BKLkpUaGejxzfFChZWX1zq
vN+fbHk+DahnXTMHRKt8FWJ77wJQBDY67mzwSoAkhHP5MGUOWBL2DTZPjYiesrkIDpaXEB0JtufX
SOoULenz6b3lu8Nf1HkLbSfGyVVpnfaP/eTNUJj2Il2Ro08/JWOmeLw3CkVF80Qvg0jrrJBdleGN
tDT7roi5YyRcVIp/Ys0XvNLOtUF0Dw/aoO7ehXfGCQnekDsSBQeZPEwOOiOAgBdRVnyM6RUlltPl
s7y8BYOvBeD4g8q6EC8DYu5r7uDxB5OYpO7VPHSaxlRz7tGnkuxCUsXVVFKXJKKjoumU1xPd0BS5
LY/XbvUqfkLz+bOMJccOICFl931PvkPh2jeYsX517MMcucvnBZDxQTZ/w6Jed9MuwSp9pVlMcRXC
R5atuO7Wm9v/oz5pyrDp+PUBan+FaobUus0QUJ9aepr2jGPHF7qf6x1VDiJZ+FstJztIETKyaE/T
scUO57ISuClBa+KRHMEtybQ9HLQaoz/HMG0D5JL09gwqgU5UlF9FaldLvTDAbjiM4eMAJ4YAjQ2x
5OPlUKGLmhBZtlMv1oLZGxO2IX6nIITykLInEGtRCLEktYkg8NiRk5qAL2wxYSOaOoFLyrFw5U20
voGNkS7dqcjVIyQd1SNVv9bnjYVtEK4uemgmBdIS2H/y0Axx0FMy9qhnwzXSuEpCq9oNQoTPwQ1w
2fzxg/FC4GGFvLHnst/N3e9vZ9z8v7dvjNlHb2XTfXEXFmC8G88C+ZxUIAJpWM3WaCUluZm7P+oJ
XQxIGB8O1mmfITzvA0n5RgvF6JUu+xnrlj18LH2r6paGOlpQuMRmNIm+nPA4TvfsW23FDp4/UMPP
q3hVRdITxASEDz4ng1tldc59bcntJ+hb1yECh32685V7Ifi5xNomnAfW4PzPzHmfJplisEiB9MGf
MDAhZwikbo3jOnkpb6/Ri6ZgeO2Ta9Up6g2fPOXXBiiAbBt0AxOMc3QNB3PH9+huaHdubIDoGqNj
mP+DSAfzePLM/S4JMfbHJsRMz3++2lqdES7L/1Yq3rAxjYJTp4EpGZFekIFZF5wFZwnbqbGEB5mp
B4WB5dKAeh6tH7/aUuDOosp0Ef0RKbG/dlP0gnzfxedxJhUnLIDDpq68R+ZgSJVG2T31hHdBeEXZ
NbJ5aLZshPQpg9KCsI98n5wgOadwARFahFYv7NmVWqR//v/JahOtlBBvdDtTOfzz5LxuOS3c/qp0
rj9/O/tQ+VVsq8Oj4dmEsBZsxU3yXKnwcGBV74DvjuekqMRnN4XbhLr6EAV911qAonAng1pioygO
LejeATmAeCFwOa1RLtns3eY7QmY5I9aO1ttVYu+VougRSDcnrgdwbKDUL6gZK4r4Lg8ro7t1RdQ3
nAa+Ux/QhVZ/YvnrIOVlsTmZNhqpZJHTbL+zoYM6c+AnM8pvS/wdZT4K8/E8t6R0BX1cuqcpvHED
ZzUkvQLBRUMDNycwubnQdr0zHi/Y1VsJFWwCiohMEMIkTfRl7P04GJB9go7NdLpuIygphIwKqoyy
TH0xfPRRjdt2UBvmJOG8IHqseOj8+HqThE72AOs6MkMD99Ao7kp/V8X988+hurLHPwwRa0JgyvEo
RZnegvvRwEjuFVZudoHBNvL+klKM7lQj23gUtZM6kPshcJ43BUNulN9+SRfkFXL0uUbQdkJ/35E0
Mcvo8Fh5ohMPWEIheiikO5pCdCvmtWAO5huUThCSWY0XGi2x16veLEsqCIwEeY5JgONGax61/J+3
mkSd5BBehegtYlOxdKm/D3UMRg3tda2Pt8JE1jXgWP4jdpgCC3rIFMAkVCWfb9olgNqwXw87KjXA
9y+BsPzh+0wo9NdCwXC3Oa2Ed0ECgQlCsAOKihVC7pwgeszT0AwI1/HC1aNZg6888A10d1iU7yBa
XovfzpbwdFjJF7Y1lhr/MLCNNw80KdaX0Iyq9N1IZy9qFhQFyl5iiDBmtUFCOoGbGlYc9d9u0Vd8
0oXyDFq5Xa5JbVB+LorPEJfm1NbTr/+P1Lvii5ml04e2I4MQpxhHzNKIeWBAdSNNkk1FrY6ayd4T
5sK6Y1vTAI3wl/dSG6WFaniY9DzJhYZgjUoDnUMhxgYGcU6lF9SXWHeFzQDWZ7GMb+9MavYqUwHG
YcSR2e3Hmx1EZva0vlldPHx1OFh8SmXKUwpYJdErFu0BQxrgQXQ9OjfcLNduw1x9uBMZVKzCNGkr
zPxB/ZEfAePx6DsAf8GKAvvdhMrqARnleE95VbwBG57WG9M7ch15dgNWg4feJd30DhIXMMvqWFWy
U7svGLUGX9zCrNU+WwXWOnHas3pML96nUKTUqKuKuB4+y2iB5ivUNDrjZpsFM4BlH/xH4yWNVgAz
LVyYTDQO+VfKODCYFJgXAVlYoSpCdpKeruFBo7FT+Auom58Qbi26X+DJuHRqvDPBULYvtqjsagYf
MGVewk1WuPxL/mFalgncsMMuvnmkXUAO6m8nMP5LbiP3GGLpP77QqyOICUsQBN9NN9I+GwSnqwDl
PrCS0NXS7NTcUiucucqcHgQoE9DuuykO6ki4eitgfB6CP1uPZOlqVQrr8VIobEasISeLB7wCtuOQ
SlA/B2Mrw8DTIQPGlPxdLWwxlxKniS8RHYbjKFg8fmpqDRK1vuNNVyzhZavlW8t74qAi26x4jlMv
vZje03dh+W/8+uWcnh72L3rFg8E/vJI2iH8DL7Ip3DBUUK+w3gre3DYoOtEsp+EQA/ybRtj0gRCb
mxP0mdLzFm32rx04LG/qAXt9ceV+aJVW5O/AfPD4cJnCe6fAH1klm2zfTfHA3V+PCTUBVMih6zF6
o7UJiQ7GJI3ZvSGUvd6GD0r3vZG9PJ5sIKoPLKoJZ2//we9wH+j0mIq/i6KU854QDvnTNZYQHzdm
NpG7oVbA091dIOaFPlP8dDieHlH6FaW136QetB8xEqEgT6Y/E/j1noprQRgr9/TsKpdzQTmj6mNU
piaYVscDNs8UDOcm8P0Cd7QnjdvLqJfkwaALpL/VNfdsKxL6hKOixC5WiwMAsRvTpDkE+QV7uH+P
NwJBGhLv/4RojPmHq1zFnzy4/qVmH8OhnollxzzvGNhl1ckjnYCRYMcbP8Yw9OhhyLAFucrfQlyS
NyS4CpHMx2WWi3M//pTUhNbFEkCOkAkSXlu6fRNAVLFTuIzZfLhS3Fad0bISP82Y/px85jyS6S9F
2l5HxKvcmK0SjmmRuqbG+8mihfAbxKdwLox4beK4VLw5OfOnoK841drIk8/x/UTNJAVr+fAagksb
anir430GpQyRPSBPOuyDtFuT2XXc/0Pwgw5VxOB00Y6D7E2vP36iWpyBnJPGXAZ2U47Y7d42ZMQD
1ZjuBlcgVLsHbKixqmZjzsd8jMqv/WEMKJ8ymaKDme/RPcdx+Eto/0PTT1Au8ZKKQuyTOEPzlM5L
CSsVPqujbONHBaCz4lK/uRTahZOn6yw4mZkty7WHrdOC44PbKpEiQrHoZjq9bkLsNz0p94NoQa69
++kUrNg+3UuxC+sPCB3nCI0k+ONCm2qSPIwiYESqawKapJSM4jGjNEdLsHhvhCXHMcQeSkVPaIkr
thdz0GZ7eHMlj/PVGzdrKXHVDkd9Sel0wReVsSYJkE8uoJ2yR+hEmqHdk/+zn1R6lhqClq1/oz8c
2M6uc8bkyGPZtW8uH7ppFhE+oauWYc4R4zSd1Vi2twSmU61ex0PrpdUNk6r60GQmjYmaHux8oHwM
Fg24WX/8s04wvQfUkvv2x8hqW832yArKBDtZf+4u842+GjKwG7Z1zfBNeNYm7jQTEISYjrZCxnf2
g5cZQgr8DpZfGvc2MiOal8KM8TGs0d6mPKJXm+POFVg0PYt7437OIgxv2u80GJiPvicRZslfP+Cd
kRdaPcPiOARevn5fWt8X2AaE4Zts6WFxqdOTbbFUw80IqVZaACAxQoLH8acFuE48oYZqotvCqUMT
I3b9Yr/NPu/BG1CxWKPkU8KqZxY7uEhWQny4fbo4WpMHHt/z1LOhSclldyxJjb60JA0buvYJKNYd
qNmm8uxTzblx/5Ydp3d+dwPgfD+mRukehGHjySwE6C7j1+Ofa0lDq6HMrmPUI1RNO+1fA0q2PPJ6
fPZeI1yLz1u18KI0bnCJshvmPj6P8qSt5cMjmHadbOV56NdV+LN+de2vBtzUSk6XuyW96azbJiBe
kovbwlmlBSZ2q5v+hck8xyeF95ILMKFKQMrqWh+iyvIoRvCjlKQdVwWvlD7dGHKqXuQ+e0j4/8ed
TROLL/fK2O0c5nx2tfY4KhlQyAxqB0BMlwdHhWHHKEob3I95nUcu0DfVXShZxxbMRBrCrWHEBhUa
4WnBJPwnpyc5SQNb7jpPhiN+zwlkrOzo9EHiWMEoQlecfIFAsbPGiyaWxFehegyG9lb/TQ3i+6wV
0cruc2XJ2EGMfIkx3ys8F2fS21ZPdGF463lRMyGglLnLnePoLHXGWOCPE52w8+GwnkEzQGS84rQI
iFGFHxDAdhuGn/4Oq8cA/SCaW4mMSN/ljM97FDMnIC8mUZQes79KZW/PswADd4bQG/Q4/YLoETqR
bAVmCzK+gnBLu2x6XASZSVt5PWh2ZuVLP+paKNsnaiQiyEAReG/NUc2oxyv8WrTDdxx6kiLPB4iS
CUaRalUX0QkfPAdThTkjz8Ic6K1WXTyFy6dqmQ6XJEizT0C/rgw6fzxs78+HKRDWzfR5tCUAfMxa
3r30a/ijPcO7oIm5oRD1+oFaxw6E97v4OG+hspHfycmSSrT/ojsT1WFpYWNvKApTcaiaiF2jiz1s
Q9+lgUsWPrWc97tAhl2uNaE3blfq9H5VHPeecfpWCQFYmGwtgDtw7vDTjobPcc4ukKoHL+3rLJVq
MPDcQi14XMaoQwWbP8I8Inr5YKzLxEWf8Ud5QDG6qDTCLyJCp1UD4Hi/zPPO5966uDJv7hsoxXSI
shI9j9LSRPiZSbBj9Ijdh8y6msvqzOxhuiqJkJZ4mXy5sjagCGGWQjZ0DtbBIY/3EY506t4S3udI
OLK1BCOLBjXZKoDH0n5nN3AI26m9BpFoHZJkQa2Bqvo4FV/a3xr68In+uo5HzFMVGv/+spaj0H3w
yxGW9JQGywG3IZK/FPYQAuO59HOP9ro23mnZs3SpPoFrTmp2Glfj5mxV22daxbpLv+0IKurPgeLA
Vnu3Bo1aRrqa9PbLFXH7lZVaITEheMr7gTU10pLoPlIWBr55FhnImjr9n47oD+7d7S6RQwzpfqeM
qZrmmjfk2nPEiCYbjTD9/cibrOzcrDHeLvhF+3y6yOAzV9XtVYjt1yg+Cusi8WjYFJpgGu0YBgha
0tfCBq74Iya5xbfKQodnZl7dWUF1VQR5nVMZMzahCIuQQ6Xu3VnDucbAZCxVkdSKyu0DxXp+m+Ru
kAEOW1kyAOcNA+Zx1+EKa2sVlx3LW+7VlQRd3xyTyiQMcVndu+3M+7XyGsE7X8EleqEVuzVFuEWW
Twp6tg1LE5+5l6I7pFvkCTT2jgNXgmp6t/YL+9eFOHKyD5r3i9Sx0HOHVdlR0GvlY9zNUrKfmGHx
vsbvjepl+Zy44/AgdpngwWerxhPlzxr2Ou6x9morArq3Jt2L7CAAC6Quhrp+013CfAFh/G8Zi5XW
wRi3vShm3hyZeWtUn49dXMOpVwaDJizvaghgfrII5F6setPNl//tAV5lLLHA/3/s9ygdWqV43AVd
NEnDPos1OJPCom1cZvNByGlE5ovBiRXVH9p1qIZ006+P8DbR71cVv3FzNdL7+Y8qYW+/BgW2FO7r
rDh1v/kPW1XcolEhPbt59J0uPJF/IruyA4MXUB2KGC5a7fpP+HCAO6U5wNQPSfXhldxwAjyz+nxk
ltI9UfKMet7nazRuGUxaiqhdxFP+Yg6h2bD9W1vHyqkDJUPDIH4dvr4oQmLRJJU49AQiIYKadWoz
Z7GGg+LpOWrkDoxt63sJz1OLuLqxuhMmpfENj2hi814xJ0zBBkT4xuPnfTgvP3w4o1t/LZfjOklZ
Mp7hlILui7MyyjG0VgOyKlx2lgIvuDnjlwxijSS1Qf48nQroY3weHoI+M5UVrJIS13c5nSctjeDs
N6lbXLyNyXk3xx0oHsaJ5oxECAeGbBKqBM4+eWTx+iFqk79CMS8zSstpi5ypqx2Ab+r8CnIByN03
Kc9h5m7sgdqS/FWU77xU/NDnmkEk/ajTbIj5VfKSqphwvNIGurIlfYIvpb4aLzOCpjRgn0gM7Pxm
FjPY7RkAaqxf3jTluOROd4s5vtXvIlhRBIiS+aInQ0hzDT64DWe8GhfwAFDGeegwJDge206BNLpz
IDW6YiWX/4pXgI/J2H63fvkS+CHuzYOaDiSUXE9UE83Zn2wY8xV5/pcorhDNpH+tQiH7UWoC+0sV
OXzTtNIlhYeK/QkAV+vlsTFLvEsL/EqgvOs/RtQQZVfOgEpMHkjLozGGqM2jvxH2moKF/ulypCAa
tTs1O1RDzDCkJlJG1yfou4FjHEnH9c2xdhblMN41VO/6W1SCzmTwBS0UZHAmY3ECFJJxZnxdGvWT
lQLZT681KVxCtVeOFKk9i50byUdvwuNMXO6u+hvPTQ21/KdaqY1jFO+pT6eh4aKJP5HDUpXnDUuD
V4D4Ztbl5zl8v0egbcSyb9rerJuZtGAUB7U65+UY3RDavOMIhrmKDU3VYpbEatSkigDr07oljd5D
9t9yALWUYq3DP7W+S1T2q0fldIskMNdccxzN8kz7HmHPSOrTflPQzfzeyaDLY7S/dgFqLrpQ+rcD
o+BS968L5/3/Xd0QvAVbQKQi0+RcVQ6zoZlIbkZWrs+W72GUqkcFaJZOOyEXhSA8cEA/yPcyTZSE
vi0R4ExiPpujQ4inLE6gGFISjBtFQdSWbcaUkj8PdNJg2dSnIRzTjMc/5mqE3l8MHj1Hrvm5JjX1
7xiWJAEL7cX7RGqH823URRLCEabOje6NLElBp8Fc7yjYCENqq53q1SJ8L1duuRYTJeASNnhovnZF
1ZtXoo2pmiQbcqPoaRnyZV4mcDNmoWSjWvlLOBRG2+QLcWMZuL+e+QbGPMwlxv68KJieRZ73XqY+
vbPKhmRCCwEiihFSIMTF5Jwmpa2MQArL6nL/j0eu7Mr01r9Qbp/UQ5GgeE4DRDvCFoYRw6Xge5TW
JmryReYT/biQw1mN0sEXlxVuKpY3juvLJW00rLGIcNKyjrLeHX1Dy0pbyiovksOJpdGaIEz4U0ca
zKEsJQ+3CFmNzNIUiOD1vFY0FWg1SEWh+8vzXPw9LJ4TPQuAk28A/o/8xZHTAgK7bJZ5k8c9HGfy
yfy7T3sHVgS3adK/0pEupCqHsy/6b2poLMlUJM7t4DDMXJHe/MEqOy4Vz7hsubGoqTMvVtHG0fze
Nb7gHIp/sKCWuPKfDRCX/as9X0nuYQt6rFB5+77B/jWzGljZRNKMR7XJO/KRoiNEY6mIYzOkzk2q
V5t1RLIpgiD8HMTwrtty3tlXUTeemMJpdwAWt/I9oNJNJfV1ahgUFn8+dbmG/akOm4caaqN0vPJm
8/Nv322mF4kCyGJOt8oMfityBnhl0g8wQdOG/AXhZIh6Hfxzb3PxAgnp+HtbmCzH29sTMvs4Rkc2
/SxIqNhvD6f+PzPoA56uNAX1jBfJzLVWQRAG7Kwb5MGFZZmTVcNf+7tlAkIMKwWKXmXAesMIdZMp
k2NFm5bU/qzgbkPa8naO/oLNZ1a5GnpYTnA0T0Vbb2YeoIDLuPGjI5Mox887tp3/s1OC27IZigM1
2wbQbmKgjWiAI2eZhJAqKc+l5Xw6O6pzAi3D0dKy5VMoQfqp73psdiUUFKHqthR7InJnlXKHssiU
qBukIGTWi2b/TOl8lrYb2M3lQC3PIT379AYZDaS8ZTRkF/zjye0/f4mmvJ6T9kHPpTxjAeZzw4Jr
q1413WfM5HqHaCoMt4cATnuEFCcy6g/sOzFrwe50em6H2Mbjy7Au/fR9SCtOMpvS4KRAGEkMP/LG
sQZ8qpGbPSWTuqsZISh1M9uz8SzmXOl5qbQUFDH6EaUO1sQp2MEhGtBEcy0lheB7dO7IR8mig92o
LHxROx6TtNmBXpUoVBWRQWqoTAM+K+Z8GJaxigsvgmvVA9f+H/GvWh/253BMjaDzCGnIAqkhOcyn
QgAQNefTDED3B29QfMNRiKVMFWzjs5ihaR/ma+QfqB9d9xqmoF6ztY3pDcob4sF2vW/leXVSG9hL
OSx3Ba8wNARFscJ+/ct0vOZ40s75UEgNnPMXgnZ6/jgywESvexzR5BMF3ys+2wlkHGWcvJX/Oe4t
lvRguVl5f448iZrkwmuAVO2HLEJJ9k+khMnQla3mAubDazDVi9dXcmSho5UHRSqQbBhSzMB4u/00
r/NGO9EN2PbEQMWLD2U0nNM0Yn/RmluP6GKLwqh2soWOSRHQ9SNDthJm9M7sCbXe3GxVKAzuLzop
7NrwjG5i2A/oiO8Hai6sM3ULZsjEHeUGD51SEC9m0i8ADyNKNHxK6kGQcEMLylpm0/htvh6hpS46
aeM/D1ddf0ijiWApFivL9h08mx74f8giKwderIquLmnruTnMihPyHXt5eFv8G+gE91gxFSTQFuv7
UZMzmZTuMIj8UaLVTRxWVTmj3PFAw1qHvGJsOPsNCBjrLu/WDCqlABTcModM09stj+LirM4dzHgX
yzyX5aNx5/PQz+Q4di939Xt3Lw9k205gQW/hitNDLPf5wHokLzQQiyK+28AVanWHeChmzSf7G5W3
LIHZxwAaaPmb3WL9wdSUAsnFwnLyP7AQTkX5l0izKHaizCwKX7KY1g8+ikVaQfkMQzeh8n+0BaaV
PO42kQgJLnSIQaVxIy8GwDJVGlbu80ikZjJgenV51ZgjpunQ1Lvl7w6KM2Z5PV0mZlsK6yz3toBG
2uwclkPhFB9qMsueJ/WrKmO9O73wWiPi508uP3hrH2pfBcPg/JZNlmnHR6MayBFBz14+wRtn29xb
I1w7JoCvfwIgic1BWxx++dg26uV+opchZk71W32dXQlkaHoL3NvB4qa06rWWMXTSHKNla6kC0pNH
ozQ58kg8sa8sXtcqyDDrl5+LLpuRO4gGoP/IwwRIOdmnrT1d0aOtE2zP3hOnrdXhx9vPyRPNoORv
hQdv8divlydcEdvLLSNFHYtLplNDVs0robglpRr+FQ5mSTSnxH9ah7vUoS470RJNgiJSFS+LKDfs
leU4I2KTX31QALwPkB/ZQYmJDY65wE5E7ML6vllUWgLh88FwGu9VLkD4cT2V6Xu+DW33b9BheWrI
RkIP2HaMxE4LOqLpYgmqzyHCZA9tdSw4nyw2EuhOzyn47bjwyo1Cftr0tnbMqPm+MKULR//PFQ9c
I+MUYxjHxOqxq1gLC5hkDoXxkxNNJaigoAWO0eQWwAV2UZASD6Mjfql1Fw+WcOrr82Q43UeT/+6E
cZ4hYQ46pmudivs9zdzY9/EmYuzMPMKUGW5I/8R2CXFXdmaZU2KkFge8imqtVI9GVUtSdcNIGlCW
EVEMcskQ4rbCU0Ty2+LYfSZ1SAMjJEOaeaJcZjzhtdRcj5CRJJnK22+WBuLf73mxhU3vFkqxJq7+
mHq4PQ1AjJBmpZ5W2ZIWN9xpT56rzi7T74FVJyF8AzSR3gC+MJXouKLyL/kmZkzUP8btMJl96yki
+8xqDSS4zvi91RN67aJIARuUIXoM96ydf9eIzFbmAhYd7ZfesWReBPuu88ImjsV0XTOdyJMhkh34
+3R2Wr7L19xRWyVuy8Ljvd7Or5Una0QQPZxY/wVo7FBrxqUHcE5RQxHrTydo9Mi5ydpQxXErNh8x
Tq5kZuRSL4sFwVOmOGaEwBYo4s7H1ejhPzoRNYc9dupn05q7uv9RXJzht2H6zQOjDgnMqcFeaN3d
ZIQUB7u7jnbHBJqK6xkL5qtY0wr2KmkpyGOLqBipSVAnCkxrI2myJfpg1SJaz3Y1wlkip7GyP0c/
WUh0pPorA+5mq6Hde+rxXPC7VmNqhh1zW3Oi3iXqTiwJvD840tLUOnPiBzLaQCmPNN/OXZPbcxWb
tOxAQZYeR/2R3+u7S0KgKgfzrLR08yyvDfU0P5M+FNwMLUTLa8AwZuZSJfCzomVvBu89WyfF1Uen
m+2L7l2SBD1UcgZN0Br13RimYI1AZZnbOI8+3zvV4mL4eFQ0Tvjf2VbU1P++UZU5xp9ARhWwJGOp
jnedO89DQ1/a8a/z/gQk5TXfiLo1A6a+GTp/CGl9gnz5aodVFCnAiiEOG1+udn/1fgwZU4leNAWC
RbsoYYULl/UYhhrTI25UjxV4tc5TDUsPszyrID70Cc/NT4OPSbSajWy14jTbAbaSs+XFp8wpfHD+
nONpog2pwj/hz3Xt10fvVjinJwFZHE1PC70YkkX+Yf4a/q01g2VGK7ghFxlVJg6tIYDuN3xsaZjr
y1W8lsTuu6kfOAPVK90260dyYcJ43QSU4qhF+MSHpSG+3+qVMuomhUzFMq7R5phUkmYUxK/dSONs
tdTOI9KNlKHPQfxHazm2QGSY5KwqYPAwyYNq1x4IwIgmU+geC9/We8uRVZIvgMx7AJ5Ccv+itCeF
tzoOS4q/RupW2MhdPb3ZmfBeOhgf2FkecR9jiCGIEevWE3Ir/FWUVrx1BxhZt+at3gQQGef7/RGT
mMmIrisXfl5LGG4JQXSYzkE23OvWwb8CD48qrGcmLMvTfmmTZ3f0xGiwd8dLfpLUeSzMttpp/sRI
o9jXk2EjiyqTODVvy8EhlPKimvEVgcTAv+xFvMcxKtkbz25auw2+M8UYAYBahMR/DwSumk7INhMC
TwwLybbJKM0+28J6r/z1Tk/RVS0YP5VD3FH/wB+Pqc/RxJAwvePcDRtJAtT+Z9mXX9NjRNwblp9d
Alp7B5Ae6rkUE//CQL72Len4uDAFeTBDKPwCnrBxFF47pkvEXFBLk9AHLkKLprLoMZChYxmz7Hop
b84L0NW2+Pw/AtiFZV9kPw1/78Z3EAl6JpE/69cfYDyT3t8yRsVYXdkEJ/Uxs1X3gTFmzC12adIh
zBUaXeNdwnogiFKEHsfmfhqEVBUakJuG6hzoKgRM8ekMSK8pkTcDDAZpzpT3U183Vweda5CMVFmk
L1mVxphZ5VFF2zI7ZGbCm1U9wy3GHQsigyM6oy9rtZ40M2rXVv3+HvTQEKUHBwsXxEJEt2v9WXAW
DXkp5fZ7JJUg7vWBrsWk/kfJT5OgmmBxPzmk5Zq4OhuCfNraamHVMHCU7i2ox5GaD58uuKZb8BPb
++3n1BtJCT3qxsXVIqjevIyfw3cJQfbT
`pragma protect end_protected
