// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
B1VpsxucnSC1PQLPN6lmFLsWUVpED5kLvB5nRARzoNHe6xQ0obqEaxckRCCI23HEkmiFMfuiHB46
YYvyDygoQ649iOet1r2LMwRzep/ACt2Hz3asQeUovB9C7aOSuwHYm8uhz6FX4pWo6HHBmbiax4rD
ielwuV+J3F7NkBzL0x6L3PGV4CpCYFokOx+04iY1YLYgzZ3Dc0sIjh6WeXIdFkm/p3OB0R5uQqa+
TABQNBU4tB0rGQtB+uMyiqJ+JhrjIWmAkSz5RKQkYQJgJ5pCG8LvXfXtQM1PrVl0FI7B3GYksl7B
feLRVgiL5OUedpHFhbrdkwePwATRYUFtlS6OkQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 16672)
br1tTHFsrbWxqnpMCbEF3Tu0EDhyc9hy69l35AznmoWGTmqn+732XCrqIgChF7BKzdyygynvPYsX
xs9/n9qJa/lxz7ZM0ZXELjfTrEic+vtfN1ReNWfO+lyJ2mBlYP9u2GJPtiy+CQFHJ7GvKJ2XQkfo
o00a7VPCgPbVjNSrpe5LZj4JvtqIKThPF7M3EmNSzp1U9wKolMIkW6wWafamSfTL+o0iX4KNnKf6
7maUvuhDINbw09Stjr1T20gLCVZaXWORq6ekZMn2qDDrnIatz76USlYGlc1tTLEO5WjTHZFLF+JV
oypD+/ACaLMFA966TEffWmdGMir0b/1JQgD+bVrLBf+e8ur/BxlQ3I1LJds5VeYq8wi16i9UC5wy
xd18vqpU1yofIh1c6gE2SGQemeow+q5URRN1jzPnFd9QwG15t0anDJ9q97kKLmnLXs4m+wWl8WYr
1PX65/X/KTeWEOzlSbhc8shS7N9sO4JBg4YFr2WsxagRxB+wLt9/e+xjOE5LxkDgVPvTPPFvSqlF
pbewXSiLd6sWdfpZaRnu+yCXHBiJRixUkHdOuhNpUSySWOrgNg7kcOijY34waja6+RuvXCygaZ57
KmDqKrgca5UaAYNGClPRvR+W+JAdRtTlkStVl+9X6gr8E+af0ak5y2SPdEH1uiGERBNYQRWszhhI
+/LV9ojxCx6Antc1qtFn0Ty/ixa/u1bUbyhcVLiATcwCevvkLcIggNOji49ePTO0H5V8iGPCGiuc
7u5nZOvWDQPkWhG32GDcpK5zqBZAod+821yMTzifiFGRX6eEm7JJJP8yLpKNlYr0Ma8lrtqLcmdx
7tYwx9cVIRVXxKdTP8aIynuHCTJ+/gcLm818a20UUknAFguBqzG71oEZQ30bR/QRFsVeZ+PS71zq
1sq1ryqVbp0P1WjfDQFxN39dwuGegWhbDL1f2ph7IBziNKp0VovpjzcJnKCnJwuGCsac8Ubz8C4+
2Jz2PGODy69LLrHJxzKJwBnEiWOoNBHPPb2VI9AbCzAF+VKdibUcmFoqfsNZRmIO1HMSBDqUC6tH
qkqiikEdmd5SfOnAIXBX5OIfsZf7rXiJgiEafZYnXq8YFe4im223FeiIIM3gF1E+wwGQvYhKK3rP
v0yFyGY/qZp6uUeUzD1vw6HTHmn8XbTcyRokRmj655dl1spIWSwIBjvQx9XXmM5NMILSgst/ejIi
ucMN/jgr48MbH3CKm+CLMCGIgI14CfzNE6VB6I1mYjjQyzVk0SmH2CVv4M9UcYP7gRt7Pw0Q+aq4
0pPUe9Tzx8epgvOVKpR/SliFICf/D2hnQTy8EEkIOtVSXIDPu58gPJwcuby/wR+mMFwUUSQAmh6/
gTWnLmC939WAgLUP3egN1EwzytVMh1pvhsd4QBwB/4CErrh40zBsl4nTa2WcsTNjEXvsukK+Y5AI
pXmecUSPd1+FQC4irBtmwj0U0ciwjOIK82u4kLj2bmtt6/Ne66Z+mw1LnybA5ToBEbgdRRH5qCYB
ED7m5pGXDYZ1WKtDxoBqcPOw/DWFXfPlJd76ddaYy5Uhdfdk35wza2gR4+fV1dLsXkSNU6UzCsP9
2JeCjK28kQiKTQl3h/xpbzuGj5XY9JUO2K9CzK+rQgGZEVdBLrPDF6XMKk9T8kGw30bqnlieIqG9
g3X4A+USmSLK7JzWRsAI/LIJZ39CS2/53/dsSGKI2abLqdUfxrhwmkNaTpycyFc41uCjG9KVa/gf
GmfHmevuRU/nsVHstZPFrDwWIuvhA8TWNeg8cEWZ9J9uoO2y6y8mGe0n7ogwiKRP6FzatPUeRWtf
8CA/v3Fkk9fMao1LO42kOq7fn0tuBLb8R0jTqhmQRgWTjRmOOZiMpOFcwrlnme7g8L+FojYr1wsG
Js3MYDBccWFXTf103ParxduIp+tC5gnEdbdnibtW5+gM5wlOxNq2rkGFpZJYIM+4SBAPj6ahKYbb
iehfxj8H3bGourQQ7MWZFGn2cHpG1Yz34Vjiuskok81BTp4k/qa0J37RC+HH6i85KNsVWK5a5sOf
qfAnF4HjBIgleXtpe3l+aY4b1MaSaFHklgx4Q4ve5N4BZ78iknOKAcgh08LdvJsjasUv4y8z8bWA
OzDiJUzhfws/+5304LrBHBD+5BJsa7JPzNaR/lVe+VhhbJueVLf+/zZ9t+6O5v+hZmtCxOb+Zb1+
cJYMIPKuut9smQqoaspi5bfma5KYmDIPGXN139d5H79DLPGTz4m5jvH1+ms5yPZqR1EwP7tUVITc
U017RkGfCswB6f9WoZB7dU2Lp9Eu1DLPxUy05Bc99AYzC5rkZoOrggQiEVIIM8hBEcg7zfz4yvK4
KXZ/BJQlqCC52SI2kmIg0PXW4FCK5UZDD2vC5pcVsKrobqEMFrmLEuBcOZ8VS/l/jLQb9+QrVQ42
IsSyMK9QsqK+iF2OfbGO59go8iqy3V6SoRbZYsQB6p8e4YduRTpSmVokiSfvOOxwWUzYep1uhzCw
/yNlMl7c3KtkhzdtxSAXmhnPxlsYhtTj0zKqcmWiIifeLvzYWK+dWyqR15+9bhxnHuFTpfRIfNUR
w4By1+m96ooovClE1ZCXUr3hfGDkhySMe7W1Nbp9BWLQ9P0yTiqD3rw4QoVhgnzJLacAFctCgyGj
6fYUuMy9uEYkhdm9R9k/EUN6ps2ygfNxkOp5m7Q7pF1uCPMtTkO9mI3aCSmugI56e6F70+kN7b1T
zpuYtCDV9P7jlLxqHhVOPNvCzQb/sI3CJoBOWqm688KLgikUMEdSpGOD+JQk435Zcq+iFOOqmVkp
ObyYuMjxSSD7Ok+wu8Gy8G7LF5NBaY+tS/ShRMyB26ZOEXKf0300XgjU1aqnw/OXChIsuuxDHB1K
z+HgyW2EvOLb5pQKnnzmIuXvza1Z5h8583Lpb1W2dSd5qsPA6NZZ1AmEtknfrjHRkERusjQVKCJ4
spYB/MnN9RTKGC6KNHCcL38h39twKUCoiCSfCN3zGfiO72HVC/7iWT9sTFDgrtDsjUw2KKQG5JVW
JHnu0xv29FyTQu4SQNTp5/wtL/QiMFhzXowJnQrQequMW7FXWFW4I+e1P+v5NQLmtCFZi1l1MPV1
ZopbuOiyUJp+iAHurY2rfZC+MqFMrf+utGQ62m9YIjV4DmVZAn0k7v1foaUAUT3U/xNrvNjIfMZq
5Hk8R2Ome/n6E48s2uLFJMvILVgqMirLEZGOhQO3Ahdolqz+VJhTFuHI1Ap7dKHwjHBIGegjpsii
I2i1wAG45PyrFYz8teXMUC3nIj824prk/cTYN5nXjFkYt3wDT+ksuchKoUgRQ9czUkcDENglrodZ
fiJoOD6fclKPnwFrt5vs9b8x2+uLSdKNGaBXgvjwwfUk1RFzb6RnNVpneF2QVcwC/HfkZVl1+uCX
MsMGb/a9tJ2tFfAAsGMO4101dAqHelrCOdvCKdKiySYXRI6KcA08r13VZjaD3VuT/+EFu8cyirRS
87VeIe1Iyis5XxOEwIiTpMT/WXE+Gq+EAhibBtK5d9YsRHDz/Y/dI6ZtusE2p00HfagXJ8Z3RneV
OXjohgGy6ynnUB0j0daIhpANmXGwEZ+jpIZu9ad2Ng5iud3XJXR/C4G+4b7KkjS1P4Fs/vTrOUvo
IloEpMKx1vAmvU86tw9i0twrz0/QTYBtDRGO2qO/hePARt+62KQusuV0hULG/vDh07Vl7rYazuN7
GoINak/YnKiky+TnFy+ym9xD011GAOxsyvV+yl/nfXvCxXR+0OdpHaYUyRfHp6rBfI7hy7sYF6Dp
8Lh7jiRJ3aejgY4fNen+y8CLRmxnp0pX/8OgBSzX4q8Lige2WC1c/TnKOFXY9weILrFmPgDInPNe
j8NfhlpJl2orZraiPI23QrX60SSCbHV2i6kwgAP1A+1h4JCz+CTxmpMXMgboscXC1gmT9aY9yj64
huT3IUlBADaZeMVVAR0Kpty+Sw+zu88IFonfvByPYTKyI2W2ByBB6F0jeHHbF87d5Y4uO9RmJ7g9
YdfVTMhnByD4vY3cMNBYI9tX4n+89A4R7hYsFNxyLsat+0vFpIqU/hkzvRBllEUMEvH9Q2qkj1Ug
Ez3tEU6t2W3qdl+wmBQo+sl6eyrzuXdGOBgGyo3sDosILYkIvCmXl/w/8FRQriAVqhM1NWkuSIHQ
P+PXLlZsTVgjvBBSQ5Pks5K5poeaDA9JVFpZpV2dPLt+8gKQReT1nd3qyqe+0sR6YJGWvAv5zad0
GKPTwxvKvUTbEe4n0VRmMoJnxC+J2YzLu6RFMUIELjS1HgkSWCybJelKwOTi1SBJIu+rENjfZ0N+
z2UUk24TiTQXfEoAvkZ+xXxSXsL6ObYABWGwD207aIaLT9GMKNtYvfi80EBmAzIfSi6mNdZSZkmd
1u2NWmQtaiVH2sQViPMnWR+As4GaKc5ctLP5K5lENpM8aqWWJwDMZ4aa2UgeWKmHBPIHYsR6l0Vy
2Wl8EfRmrXc7u0fdXuxPX+8sjT2HxjVFLXAWHi7c25FE3X35nITIObDfsCbizhAplqZJ2b12UgH1
xUCfFDQD2aF2xKFnci/I95FUqgMpIb9ZQQc0L1mdpo7kVG5pZI0r+ITpNJaa+2K6NOhOE0KZtXFK
QcSTZCyiXafitdGYtfMcx1v5Ru4UuzoFcabRdCc01Yve+PqV/RCGr0UPxPISWq01ujucX4TyQylh
34rsWjBsPeGBTNOWxK/bfZ6Yy9zxhlChkIzMfQvM7br8GQYNSV3RzSW0/NgE4yOpzW/vP1FalIkG
tu25yQJJX3zNzHFLDWsJSH9EZ39ziR1905aG619tUU9XACd719JidkZnOOIIxikPhmcjAxDwQgsY
WGOY+RcErD3c7ygIP/0DbQyGe481zLG7fMgP81pYU9AdoPG3+wmw8u76mgpV61yYQrvhHCTN19A7
/4sHlybbZQSbqjV04O9XJoBKKkXtKG7Jwk8Nrlxuz4b/4l0aqAM7fCprANCcJLpfsTU/ffTX0+s1
lbdyrDWOKer+CZ8K2jonWbDo7/NUjzH1uVj1wdTDBL2+uuNfMN1OS6IPEG0G0OMgqTMicvK0EmDC
0Thp6RPiVe2SMu/yUw8WyO3xJ897ars1QlwFY5zLNUwIHTvdmg8qngHwZDfLUOQQDNSH6V/r9hQR
oD4wmspESSqTUGDgrqfc1V/QWGrjO6xA2vX3pmy55zPTckU5g0ZxInVpzG3Jg3mspthsFdS77MoR
9H3LBUB4B2xOzj5GAjaaQNFLTdSgvxjKj4GRp8ct3WLWq8SPNTLNzQb8s0hfaf0q4bm72ZVMur8g
xvEAXpb2GWj7mt1YQxJGEUsgS0x4CQs+h40pRGb7pzqqJo8yt2U9ypTAwBrEs8+nj1yvCGdizXM1
05yYg2RlodGIVXk7H4GC+QeVMSpmKZopGA0MRuOPkeBtZp3AecY+xalg+gbrekeaK8FtPb+N8Yij
iJ8yT0g38kXF4mrqnGyordNV9T4RXLr0QTqQ2UTp6JWUwtPBGX+/ApiZ7kVFf2+iI7mozH9p7ZdJ
jwOQkL0J5ErLSEk7Q4X31GtQXy2I25bL+yALYCsNHSIqxKJUyYqX1k4Je5qraHlC86xlp87MkdG3
Y1YhhPufMOn3R84br++US5ulQ72LwK3niyOn78hRDq5vBlfAeNQdJS0xOg17M/JcXcub/UFi2QNm
pewTjU438rdlhmQLU5mjirCknnv4WW9/j0fmy0/Q2o94PiIAAiBcYopPDb4OfLAVtP6vy8QLYYtS
PFFwCshNHw96BY/o8s+MKQGkTqMVKKwVcjeYX976084G4MJ/MjV0bszu32DAm6nirralvcTTUxJ8
M0+sjTANKu4Cwxzbavwzfc4HJdyQx4GJBKxxzlzVblJg8qIf1FwY9tjorsCcTSeNxRIg5Sp7lHIA
YBSuc9uVHFF3JYyNQCfJ5tad+P+TJBpjmQ4alth5HjOLF2vfwzarHyddfLGrSgswDXF0FUP9HBLW
Ds9vuwpHXIPHvU/gCDNiA22UDOgmRoMpkXu4/w0v/DvdCrVljJezZDhZEEGZePvX6l4HxYIFLz1j
sWgFxV5g98YOfyrtitjIW3S8W+8tHerAGTPAe22jlMnXh5I3ugGdG4sbnCgJLDa23okXAx1DeWWn
7nmZpbvmHMR4MiaqLuEXT20yav9+EcC3M3h49CIboxVyv3BghRmHaCCgEuZzJ/AzlHVRqCbwsL4L
XaORtYfvIlV5OV3yA1lgOK4LeL/eQAQbJ4pzOK8cspGQUMvoUAm7Ph892/mReNsmwxfOiYSFU396
4rwGEmFLzXa/CPDmfTedYqkzGS4vFxCDhh+D706MQWaaSvfuYF2evKjiO5NbR6uY98q2+PHKl1rW
WYcvp3GphtGP/dPRe+yaJaqqMdS0mkTeMt2ipezfQs/FULWmWVSkneFwHnSj0wkWT61aRzqfzKvQ
vRRPQtl2aIEwH38mfiRLyEd4E102oR29d8czjAn08qQjqXtB6tlJA5HnlCjFOEnHPh0Wfuo307yZ
vZP9h511t7B2DU4rQC5G+c/eaf9NmdQwBc24dAbVqoquMlFlN9ODyf+JTBiKEcXoUf5ZXbTGOBEr
HMAv4lNA3IvCdZ+dMpV60QXzllwweDjcvbwPjlSIv/RCmSjT6hQC9ap+JHKWr1QSiMwwldu+LDoQ
Hm1CNggrEzVljp7vFwPFoucSAlD8BLWiTUd2sSmYEwyus7ubim2CSjAFFI3Zf34Bu8Dm8sYs9w2R
PqMkZBnizbCevnsfPYpFGNxiYaMT3c27ZzINIMgUvcDQCeyKTO+Im58KHyo6txRZ9CTXiPj0rezB
LmpV7asw3oq0uxkHtcert8+ZQ/9xUn1fjfNQF532sQpvUDaueHVUqrhYBAx3SGDJ1z4TUno/DajX
V+25327HTlLxBGKG51ItVnBlOhsKeLuFw1RLywCXkJReYx56Qq3QOnPQPZ4+j83JxhrRbBrIsL4V
3QFc0d3nqPoDK/UXU/ia4lxlsDSGAlogQK8D/Y31Sv7OdSYj/uUiSv/ShUKXoDYkqXWry4eo0gG3
+TyRnGvbdkCGIEyvUwYerArQQYID4QorkJy4EJIR6eKiUYRAPL4T3qfh5cnJ/8lOvbfCPmPn2kuH
bUap9a1ShUVHXc2sp425zh4bMDSFYJ7QtdKOXU9f68SEb6benklYhTRSNaMWGZ6jh5OFCo1YmaoQ
Jpje/oc9y/R5n9sDD31Sy+K0TDTOdiYouegkY77i1fuDOEGhRpGC2JGXURJO7/ErXxf26/QQdlfd
zv4syN821yOKqqDuR87xQLokCVdGcdHHaXsO+HZDcnpvphz3Uxg3xqlfrlSEJpEJeHan0bez5Gfy
B1slRtMhhVOahnj2zvDsl77PPFCYbmqAzk1XXzcdTnsvNVd88NLC5wMKInrhFNdDnSNb1MGRueAy
tOpqvd0iG5ssugRr+A7HSnik338OogmqkJxXqzbDH877DjwvkXIecuPojvXC1z+SMZQSIJG1pkKo
X7n+h01BrpPBjlSzLI9ftE0qoXUBGgKR34KR5LYmM+NQuAEH/vK2GmWJ9qZ+6WoPjN6EbnLhQmm8
TIZsR7RvLEAMrLpfzjRPrEeqp+o5UL+dL7IUfWhjvPV7ZLoapGSyzQeXKudpR1rkTmI6DMGNn7VE
+P3lJMo1Inj1EzGJk0FJY5SUS0NH2L8J42C6hjhqHInWovWl3MLYVnPHaf0Iiz/bMP8NzyVHpnwd
bqP6cTOqi4OITPTDVnX4PGHfnwA/4foK0GpL0WQbsX0JpDjZ36D/mxyxnbz9VietM5ri0orhUS0U
aj8nYH45e+1TEpD9CDnfZUWFdAhou/eawpg7OzhQY702JqNNE9qbm2gjqaAKuuwjRtI5OSYYRc1o
eLKN/MikkA5FtnEmPKgjkJO86OvQPW1NwKxi65++6BNwya8anw/Sb6IdDQbX8/o9VvyGvqjxljxp
cio9KwAoyFVqZHBZk6+rPjA4Pry8KP+MSknVlfnLIDxX4FJ2x2ZqBmMdwzkqfb6SfnK+VOltnZRc
mZ69vOwwRIZ4aCz6k2UbUJYPXmBeo0M5eNAa23bfxLiWoZLJXr4sVwOQnt/GYLs07iel2laF2kql
+Fct3cD+xcFmuiqJuJiQzgXj8Dx/VrFHsoQ0dCYsSBFfVTlFe8cuC9n1WU9617H5AutrTndimdi4
ExAFvCVw8zQbA70IZdjrw9mS/Ha+MjAun9JBhFVQa8RnKWDByM7BToSzbnqEoseBEWM9WH2gekre
y1+BvUcXC/oLHnfQ88K96lSOMnfR2lVEMMD9upFaiGecZFyWDJjrYsA4jTOUhzhgoJzIRyl28dgh
pMVVuF6zsNXx/Gmo2kwhmi6QDsX0UNPaGkXp0WaXtRxHNmRWniC76MBzvmJX1UpUWcQ0LFhtLtmF
esMy4mjWE/VkwRRKtN/zuls2z4OvkiV1l9+upgBBPI3VhDGkkZyvb7zcUBNWjHCAvcAcdcSiCljK
sp4m86Ki9PwaSwjN6Hhzye8NAh8mTB4rVGXJcM7EOsA3XqFu+t5FrpV+5jl5AtvOXd21HGdM8n2+
iK60z+uIuaiV242Dnph/idsa5GKGlFhfD7acCj77KdEXVEB/Y/Xdepz92kkZxNlAPIegwG57tjzQ
FeHvz0Z6etBO2tuF5QITdK4m5Ma9ghDQ+/0minWm3jXDxOWUhEEmxgusizb2UON14YiCwFZ6VwIV
OQR/F3zAPbNi5p43Tf7aIZuqtbSJCseJ7c4hJix3OwsTtpbGW9rSQsaH4mWeMorDrTF0TFlqpbUM
gOqUWmQLbCOFrYXwtdDN8ot/yWQBCik4Q1vpXlifcPMh0LaLkwP3oofSrx0YjqIz32N/ae1uVxC7
mYnfR7P6isip+o1frQ0ICi3g77RT4BgxU/Y2PA2y8i2m+fARnENDJkgRfctfLadFebhLeoxuqQSB
AIr2wMJLiw25zuxZIPaM/UqwpeFn3kecFt/I+F96MM5zBvGNTVJ2nPpEWhNrlNOFhhwpsfDQVUnH
zpyok5a0zh/OFn+zfESc1ODY6VQSSRt1Z6o+nSXt2LR8AvnJRZLFzKjn1rBrAjjXp+f1Z6uHDF6X
n+OFQvfRc/l2cT1h57oUu4rttJxq/DeNWFH/AtGxmzRi8qHpSXwqmrtlzVmq8uw/xbTnx17cSMA2
IINkNAdT/UIQDDxziaPlacjLkJFuIRN1uPD69CUD28pgPpIk5WxG5BAOYb5jk7K4w8zwrhJh/dUw
UYF56FNp8CJL3wMInLbKJ/q1ulqxL9acAGLSqN/BliBZs4vYslh6XORrivLCsanQG/PS5U+bCr58
TFHWWl7qP09flTIVAozuAwwo+1glFl6gikVaL09C5w5ywiRpY75T33Zvlvrs1jzqIxmjWQMUGAMK
pm33kyy3jSsw8xwzlVGKjOGEbfhOg6m15zZXwPShNS1kc/yFoRQeP5UQnGAF/pVapi/aRrDr4j4T
CO9LBwBWP2lGlZHwX1egUcAjK5Wf8w8yM56F2rbV24UKycDbpQUcJOvtq7zNfHGAaQjOM/o86GK4
q8x/QF6LiAxsysQ1wD53b9hHCSO+ZI4ocb8Sj9BkxPEKuit8ae84bAWdI9XxjX2V6oxlE9DqzZ94
PAUgYSfYB8uNLqyKosAWeqSmzoP8GhaX+yCot6EbVpvu+ECWtAfLBq5DubczBnmwMW8yll1fxRk1
PubPxhZynDd2l2XFGmJ90ACogkSUKv9QJKl2F5STCEFkQaQ3K2WwqsuBHWgL+/vVvOpz9ZyLBDnq
+eS5icUjokMUpmMvEw5Si/xGzNg164PX+LLVQSoCtiJ8xGq0KLXw2U6BtwqRToD7WOchapj9e6v5
AprmcPU1ZYsA447KWWr+G+xoZeLjotduY0YV1EU8Z07VYjplo3AiK5/M3iOdEaj9+5M3axBJFt7e
851wdtoBFJ7+w9ePnBA08Km34uhXS4M6nut8D9dQoEjh13xUzETkuQAUTdivqR56eiJeI/SdlIfE
LvfUq/niX+B3Un+aOw2OtvxRb3eabSRqVsMqBAQE1/aDQOoX13MpsBIn5+kwttCs1mTLFY6V5Gzi
7tXi2yTZ0Laj4Uy02lTjV74axD4nsNZu6xOb9cX2k71f51oXRmYyhiJDcG8/C1MlnaaeGdYXY2dM
dA42Az2miLn0qMfvuRGEwHQtKzBZeagn/xyI8l6cFKgXAUodHvHzoBPWBqsLySbHiomNPYpRskKD
HyXIkSiEjXc496s6cJJbyOh9Dxgb5TradqATWHy2PEh4LbrCicNTgBhPOpJdqJdAa+SJYxrOBgQH
jSM9Qc8lTa8nfG959s5Q/CA8gLHbK1N5pqHTuzIsE0/anCYp3jTaOusVX0c/xuuzPXhR7lv5B3F1
1A9oVL/viKo/uwE8fEt/zHNiH4ol+j7+5s98It++KsRv/nKH/+FdvGbhn0hL4vLvO9ftBZOmBHNp
dy/B+GR2Zw3nnbv9S8LCv/OEbJR+3ZgViuKqIhI92PlPoHJEO/qvp8up9T1DL2EO2ZnWKwcPC6Rr
WqOC67ZNPLvSprwe/iYuOdeC0+qJ882sHMG1iAI4H1RuOQaOf1KNcI2tQQ31iEh2f1giYXz+ctBP
+6XsJqy6+3Q412UVjckY/z39qiN2TMItlfCJgl+3L21OOI0k1+8QI0Gy1h9u0SgqE6WwJqu3dBV4
xXpnCkr3TmBy0DXQ3+zLuwBfqprMxs/rhn9SYt19pZQ/thtmCE6yfgU6h6EByhlKI1npaVOo4MBD
eTMbfy6/XJQRzWvetdFJQwopQLXfnJMCblyssXsjcnqPvSZZJUc9KEL6oACSn3gYLToNswWNbBZZ
x3U8Pr6bnocg9Hdckkt1nqKjPqAxz19hWINaYhqnG+I+4PCScN6QKDNCaAMo0GkSOlIUcwDNdfNR
CVA6cO4ODmJmxGadweGzs4pm2kEYIiOWvc98NML5DSJRKVRzsmOWue1KPaiJ6uE2NUXZMvr6nS6q
D2/nvlBer6iewIbGteFeu3i9FjzGxEdluHo5SzSZVxqVwtzOqv7K+xfMh+5Vrc5HwMOxVxOs+HRf
C90ishSvfGgL/TTHuQh++Cae8TuuopD1v4ZW0maiNW7rQVLwFztD/JA6dK6QG7Dd8WSwtQFytSPQ
MLg53czpj+Ips2k0HMS18A7h8JRoLRW8yMmDxQOWCZAytZW7dwMIgJqhRw8jVooknI1O/XuCjT+T
BEFC0fIw2cJm+Uz6krhdowcMBGYIQpG3psIXKOnUjbPrJMytTd2wZNQ7akRXzvxKe118VIN+TLYX
iBPsMfV+1sbsOG/FvH2ehZu4pFhZbDVKi03OCu3WA3petSwn8FzfsOwOI9LfqH9dtJI2tiQKgzJL
S7r9/+6rlWK2j1qtgGUjgh0djstxsECl3KkWx2YrjnBQw9MYsXMnKaHE0sxWFU5Imj4OiUDn0gbS
L9k6ApXuZ9O862qnF7wwtCgTSLanZA/wMOCl8sxtYhxAEXOD5S93w45613cy5GklhomwBxzzEXrw
7eVYO9OSmGFoMF8GqEmI/018zCe8rFxvz7FPdnOrOEVrOnheSBQ4psBE/saiuIsWANdiBm8vKR55
HV0lfDgTMfx2xnXeHKRHSSarLAsrzGsDotyNPSIHjSQbjY/UZwT9XoUIOLIIcLq3OMc8dWJ0hFaX
Nzzz5nMIgYMLvfTRvTULvo0PPlaqGXggCs3VxrVPq3GLSubR4EqiI9/+Jo83M4DWo3kJ9RnJd23E
r7DZEmJ/0y2MBZLqDQXy1Y0C2tTaBLE3rZHmqqrXVC2VBtIs3hWRwbGijs3i3nKsWlMXMEPYIkeP
JtGkarukSEn1MGxsExaq9IVAov+/daJgm7nICQepzWqBQUF2balgEWHy8jMaToVa/xhe6QGTj/F3
2QCDu5zo49C5wxhOQpejoeOpkyuSidAC/ts4yYOa5lv3jQWxaPd/vCEITl9RxW0/nJEgTqu7TAtt
V/zQ2TbxGgNrFSZKlH43Dvz0zfGJLoKQgP1Xlw98pZnBe9rFJ9mb6gsfK2Yz7BXVxZ+xWtKc4831
g70QolDvLP4IPgol9QMNdd+Khy7KQCgnjVTlrAfqvO8a+8xHQFngy2ciHbhEm78YTq8t9sYUI/5J
+kh48dRdLY8NWo+CG7+Q7Xc+5Ct/up2Uj/dNJuPLtXMcUxigXFQkmFeZlmipsP8KjQg7WhI4PHzV
5bcWLdsI1xJ6JvvhPt0J4A8kC2Vx4ZPe+mvpA+xpcO3C59YmTB382xsI+E3fG+11eh1b4kJbmTOx
8gNooN4cj0Texn1HSUGN8Q1m9F6EOShm1QdrvDx+IF9wo5kzweHCtVs3MVa8AnpH2uLwr9HuQwkR
dn6ZEdliDP67GG2Lz5DFg4WqQFlM6zbZjha0TMjZ8WgL6e5cq/XW0XwOFmTwFlb1r9JKk10iACZn
eED8b9ziP5q/75k3q8oodo+v/uZlv2Pe7b4RjCvKqObK75OKoYDVnWDcIRsk5AW0muTukv8CXd8V
WxuCWsVd2gvrrxSlTkvfiuTiNv37xKwijkcD1j9PXpxgoSivM1aAHgqnBdj5ipCFAid2neowseXA
vYq8N72gxHE2txNpHaE8jhMLyjZm4/aURbjR8h94kcWxE6/7U99s7bT4PrdWYhK4xtgILfUyybZQ
eWvUJ24VMwrHNConwlBvqi0kBidEHEkTAurHE+o+XHmJ7fak/dfyQl7xkn99uihvGrM/w8ROPh8n
Hh/UereJzphiBE+Qx/RSY45SsE4ktRqKEkmfCh4CFLLM2animBpFpDLCEA+znJ756tPUNz6TUSlu
fgIsVmo+iMWHetGHBClU530UIxGUFr1L+BjD7kI0SYxnaTF6BSmmaKhlwW2rZM5ssXJpJMLIQgCg
sd+d0tB1n8PUeI4rZpEtC3kcy+tvG0LTy/PEYBKyw8laBFwwNM0bTGLuaL7VN3HaYQZQScgydAz5
dlJyzTUwVa5rqtbpczNuU1UVEWmCq2jMs7dgaczvHt8ikAKjX75dPro3gFaiw4iyZ6ywU1DOkVd3
PejTIat2SMSCG05O4I7LWs9M9CiPscWdeQtr6OrzWmF2CNHuRfEyPenVd5cU5ZGJBgQDPvh9jMxQ
7hK9S1JE/QoqTPe0rzNe7DIRuNz3LZsUL5761Dc0j7hOmqegZJZXSTH135tPnGVtn0i+jNRgJ1z1
rTe+h9pfirNIVeZNl/37dD98D9c5aMT0LCJyo0cH+sQqk1vVybsOwTmRTH/0A93q5mX/SM/5nR1y
GC8czGOMNQ4sQFdjnUCfb3Rit82JvkKKZMvlzUfALIaMAm2XXhXRnkRJ89pCwobi8M5f/HeQP46m
8nMpnYzmKCQTA3FXGHHoppX/SlIkmVsmxGEIt9BrsuCLDYh3piAAh87NTe9PIckjpds9T98xcdlk
mW5rRIpgdLqxBtGk6BxtdDdKcS+3B4qltzdWR775HPDDwk+xEpSL8+KO267MDrArigeCl6SySqaz
CnO6ENOgP/Yz3m0kURn9HUv2kneBUkeJWjLNLqEySnoS03I/8LWFb2PCsbldypOsh4V3f2hsc0KB
ITd6SiCyg65gVUhusliMcOIgqP4HellKn2LoBh+jwzor/N7jyg0QhWC2RzeiFhTDjYSTBze1+06v
t6qPR0EqYAV1HGwEEHyLARPnYDUndRkZrHRXiDFtqk9CM+LjxsoPYpkXhkp2peu5uYRxR0soMRc3
bHwiENcVC8Axn/dQGPcKeQT7ykrEpHiFAhuxOKHZlusc+crOvU8C0pIgbFlNUCmZVqj2X9VjRPCr
joiVGEVKa9CnFwta/XHb/y2spe4tRncaJB4kYsuEhkpjAS3NYB87yYiQq6z5SUa+GRtzCTd/L1cF
HPDbC1Jhv26RZgx5rK6irnJsCBJklDHssIeJXRNtWAcx09iqpYyOc54h0SanXP+qKsUHZQQMcOQN
tb04awmthPbhVHaTIMWAlaIW7yRNeXrGiC8qdihimWT6lzl8KlaJpptP0p2/iMCkPLzSBK8SmGLJ
tUZHmA0nFTNaLw9wt2T2YlFCPp1un6X/0WFoO5JViM0vUcKpzYZ7KDd2rKVFhhJqLsINjbJW90E6
hDmE588GolHjc+xHeuXrjYO8B1/ZqkwWaHUXD9Ra2fHFR7HBjBQpTEicTTI3PouAmImhNpIBO6s8
FNai7cMHkO4DsGpHL+tBITOWVZTevKN+9GWLKdMHj87YnhwZuNjYlxRiKS3cn8FWK2HKDIDaYhKp
QTjYkHVbp1zMrZFHsr9oLc7SWG3o1XMLxsH2aJ2A6k79uTil6qO0N2GXzjn4ZT28Yi+m7G99cfEL
6WK/RVf3pwEIIJS98ZNodmaid7anHAxU8+ZETTJyMjPBEy8EBRzyoBa/tHAyzUZrFlx05iQSF57j
7cnhfg71YCvOIPHj7j/3yoklx2OzVd8Oh1ibsk3K2871f6Rhd9Oa31nIr5SByGIN38XaZoy1DhEh
UIiFz/X9awpdnJXHKSLShOgbWuAfcEF86HbxfKIjMLW+5wJ60fNtU3ek9sI9I+FMWU74GQ0gLrg1
y0cCOrdl2btXS5HuAVd/b2+VbBhbHgmy00kD8Qfv1oQ2NXanlDV4ZRcn3XqBjNQ77zrs7pSFhDc1
Eo+IhUefS2NXErPP14v/xtqlo3yDobAD3UQuNQhCIPEcrjpn/WCCsVvigBY2+uXevXzG3qb4Zczx
27QB90FAzTfTmjoyw7F/rEvELhuUboVKmp6+AVIKufq26qGz7dzfrDR+8YxfQVMaKiP6Ccp0b+RL
LuC/w/tSuogOVd/xaLqJV+ggVnc//Nh0ar78/746ftsNUX1MNMf7bd014JK+xV9gPWHp+1NWH/4s
Krhhs9w1SOjzu52rnHYVcT7aJVSQjY5a/jc4H7bAKsp3NsfZWEEZsQApyf6wpZbvvi1tM/WhLuA9
RA8+HnpjacOwZGwbPnH31s7i+Dno3txB58FtkMX0Dk8jq3c4xpGJkXYw4iwKMSptkE8/xfy6EOhz
mMRWR0EHSqKdQBMuk84NaflHJWrUtGaTG2V+D8XtJJDgpSo9PNr+VdlvYwLz5M2xnUzdj2wWGvEP
SdFzYtOEdgRhGcPs03b/9ok3TFqS2Mu0ZOZ4uNnqACxi5O16f76qgYBLKROPdPK0XsmPhczEPrSd
qlIS6NUAKgr8QKNRhC+b461xz42KUpJLHg3td3GhqbyR5G69aT7rURS9ZrEqNkucSxfeS7/GBIqe
uzEPnseFRJRDet/pL+sP9rrntWE0qIUKmrEiqFaJfPjxatx1BqAZMJ4yW2scshvEUfaTNlM58PSn
/xx1Q4jzFkEHu9Kl/UyooAE/JvRtNK6Rf0IfHFFP995FhVJeavIUdWkyyxiwRzA8Cm5ry6P0N169
Y5lqtHAIdZ74D2WHkqWJlSF4A+GoxLYWz5VtNVMrTEJK5eFu9xcjTtJiLf0JkVyf979Tpwxk5364
eJCNaJ8RcXT4nxaxw3wKTNwUEyfUWXUBcarFmSn9v974W7bKOm00vF8Pr1B4B6XrBvqGfZF/QG9f
Q0txoRyIr2jxpGHRqs1hJETJ9+mgAff5SX7xBP7/S5otVJ3rDV8FiHGmDyTvotgeHuIENfp7aUc9
rKKQN5n2UtzZdGKzzOrLy+Axog4SvJI+5RUkY9scqfT5HujkCyd8sSFcjSjQ6O+QxdiHOaCAm8Fc
WnmYrsyBO6GFGFuVVbhTsNlHg/BUpmEbVsiiR5cVJjuPYCOtrz7Nba40N0+6IAG51wxOehYY/CuT
Hber1LWgPptMDd9VBp2qKNuA/fxXUVD29bUIB54H1KuXP+dt0iniMiPfE3lZSn0uVdoZn9c8PabC
W2yYLMiJLJuWgY3Pp/8AFgxsk++WX1gX604OsV+pbMT1oWbzrSIsCZaqOCbGYGCS3sIn0TYZ4qih
ss4tHuzU5R2Tl+v16nE2TimgR5xcsmwsQk3d7avoAZxlOSLDRLWvA+jIjkFTgLFtGEy/C+k1JvIh
33KG9Hb7TPuimRxWqSPFmkdhjMaUvbM4x8XpOlj7YDP+CTwZ/Orh8qUi6tTCVQWZfvXLACvSdMvQ
uEXhn9QyGGkz9cGkp8XAOK/BYfLKWXRlslrXP+L3yAtZvkMscMXdZyKN7X4Cqsv53lk/zkm1dY8K
aOoyA77cycIF9sAqVqdyhZroSI3l5hfei+CeBZRaSzdn+ZH7+JMab96cT0VZQvuIurH909GjpWE6
JKS/sqLqtDKg+502dnW11prLZmh6Xk4UKLxlrPUbTt9lZw33MZXkebqt4DcWO+zEJ6+whaoTVdRo
v9WQzOhycb3qn1QQRpU3U0pMSrgAotkrzDRdXNzuIkiQNApQFekx+3VDFUyKQ5R27WuMyO5Wf3mx
WgTCPIkcof+IL9+DDWmsnCohKum/2zhTdAjar+sQjp+TbtSpLfH5CJ2YZlDDNIO3kaUivC1irngU
rlghPn7+FLm6+9aOtvH1WoXuD00hxfHHsN8QVv+50AUi0D0pSMD0EPJcxY6TWVgpRzKoCXdKY+AD
IR1/nV8Hy3c43p2v5iU68o6JGr3gdurd04o66P6F4fXgZGpQH68lR9logZygn1ABBVtkm2OAs05x
JdGKurpOmfjwUIgWX8HkCQe1P24v7ZAFMrYf/f2+WK2w5Ss/9ROMtGFNvsxLi81G2TugkaeTV0vH
RcnjONF+eOmAuWWPhU9S3ZGixjYRPRscNoQ+bXCJrrfhoWns/tT2bGcCnMIEBAG4ITNJY3rfs5R3
f9iqiUGsDcFMhKv0J9kKCR1LyQq6aT6daY3KumgZmxGlaQF8PZW/eeZD2+ANTRuRLJ36exd9GAiM
K9P0sd05UZxIk32PBa7MdGaBdpkewjLAPl+YzsVHbcnmYxB4dSIiYvtV3TF4hYyNtgAGSWbCTy4Y
M+3Q+XHLe+UmezVxMfRlCzwq1w0YuXjcYrIQH9USjfAhURVa21rXEc/EARkJKErf/+5RjCePEuCK
7bHByTod6P6aRPiK7WZUMp7RJ60MQBCSjJCbQ52xln+9guFDvDeYrGnkhqQYYv5xcsxcxNhzeenj
TGNyTXJ45ae3UUyi32UzDiHE1P3cws6t4VbWtYsi0+0VO8TJJZZ6uiaHJCiO+jcuD9WoDrEb3nSk
WtZgxfuNA8T0ywD8cTLo/9/K27iwIZyegLOFPyNbMX7HQI6TpQJVUiPDWCNM/HAXoSzCJU+G+YhY
xeEokcYpC4zLhAkmF7HjD+0W4dRCEAs+Eq7VNJGdvVdmgto81PupJOt4+x/MRRKMoTmY2R0B1Plh
CdWdSU6gouNc95pZ+kFjbz+AUrX1ZxsqiBXownIeMoWVH2kP5jRQdfXS0Y1VVjCPrxPniZJpCIhq
51WOMyChmm/cG7hCif9zWl0Vl6htBhi1z/sxpJ7UDS1V0brrxJjIskk1DsupCqRpK8mjOTnXNl5L
ldliKfIkjOwI8pS4U6e+BRH4PPbFaqPdIsnQ8lVRvTk/1Y/54xzO9Eax/2g6hdo4utXeQkwKOh6j
M/k3P/egSjCIARPmGdBX5A8H9ZEvd8K21PUuyn/jjiBQDMlY0CnMyLqZ5BJf4MZR1qW6A3mfE7Dn
SYbOB8+rljLb6RF5UBTV6WWK9hy/QFBNFOcuUC+9841og0PJJDUhu/YVRpbqL1z7gicv6uiqLZlj
IIozEWeC7n9y8J59B2p0bxG8ZpfdeCZ8rID21Bs4dh/iw85psa3DJol5ImIkyZ4PuOt0OY2K/4RG
gMTRSqUHXOvmrc1j//ewq+GlmUbEYqbom1jbHpIR1UXedIk8r6mB1r9N/Ab57jDNqtX1pTPJb3IW
yLUHRPgyBgyzlHiSqNDVay/rZpeNQH4r4QKvSWsMH31bO/xL0b4nT036OPwRPzXj4JjcdW5Eu++/
sOu4FzOZD/7xPzsDn7yl11caEuHcvzEYKFtx7dVSjHH/PIvSktLtob4mhs1DMR6sB/E5UYZPQNxX
WmPcvr+JBOChiHYcKaTe6SgHR3eoO6g2udZ6mubY9IiTEVyCWr/F/CMCA373gANlLzuSgL/3jyMj
1FUau+s3oWvTXUFmAf7sVxfndFeCWO2zqaboG6iey4bQ+mZ8Rtvsel45ZLVEBBanFfZ/7L0voEje
TA04M54lOw1c7/dFK4YXztuajEl9kRNqZldBL4pCHZB+7Ih7gYBna+CPlB6xhxdpl+MffGz+wqL4
JbUdMEYmSwQIDVB69Tz/mE2z/AMS8qz0gQRiwM9cNAo6Ddo45OOkDpDRcL6m3nR2WiGxM5XITyWz
C1hMO5rjS/DMiV5I98AK3TmmEnFZ6RsB4R5gr9TTjpCUOmFsVMPa8azrxXG16INXwD1UmVehcFqM
kgPamEpKNpatuLs1xpTgdfIHeKEdLGJnB/RAS/LJaBppT+IGImQQjh6wfyEXrmgO19lT0fuZ7sBk
5tOpnJaKR/kGoe9ZWazwLLphbQ0geeIlpxyDagWqqh8fyKOMcKI7r2tK//E8sjELB/Jtiiz1mKJq
AYY2eCxKjgmppiP4a9o7aon5M/Rj20wrSgNfpLuWFpjvckXUvyKaXetwBBe7A9+oDSktshv+pQFF
1NtoQL02D7qeQMAi92/7oLb1GAPYJEkpuKMIo7mx1/3+6ATsuFKO5sM2uKpRFEP8sm1zDSOTbxgY
1Hv/i0CuvvrI2aB0EBiyw1k9L/7W57IOXMv9H9uaRZFY2lp0/AxyDAY1YF1utxWVm15cMO6UmTNW
XzM5PzWIE1vvLFMFQfRQGXSaJbn2fbwt0d8R5gGtu5j2I7JrLoqaYrlKuHMf0s9pKqF52Heystie
r2UyQBxQYmPCh+zzDhIvMazpbiuDZ03+MBpG+ls90vW+o3iT3vbxRDlahIg51pROI5qMXvBJ03S6
fE0tKY8jAp6Lyz6MMRIV9fqq0ellQsyjjs4iQ0YnnPjpR2NuKvRT5awF5Jmjv0D3P5IZ8f4Ql+r4
tCf4xF9IONRDBR1P/Qgh1ChCAlAWAIGzgKbQFbywRI77fmdBMKlCybYOrDFJwY7Y5OAQei/1W8SB
pvTDtZvRSAKbI4zQ7xd6Y+zcKZpemV0Gz/Js2/gVYEoPUXRTOsmZSqwcyqHXq0PGFEP7myfGsdXH
ASZ2ErPTGbEmPLtGW1myEx54G4G65NhRB4xmWPRjve5nM6XTMoEIMyqskwudHCoBRr+FTUadvwbB
0a4k6L0G9I22qaafE/8dpO7/TG4JpIjm/RjQHc19alRNSLdabBgvP///FTXB2iCMxhCk6VgHMDCT
JoMxdttxQQsONwxqrSv517hdz1OAJNyOr9oaUxz61RVHQI1pNMOA+FcL5Upw7ZXOcVv1Rlpp6rAg
yHqIhuzfFf1gd4XoXEIF7Y9uMzFgSogKYSgzjOAH8LXJbCHqUpbIziFH00N3Wg2BtTw3LYU6WNRy
Wv92+dRfYUhjO44VdZv/+1mbLmGLdwbCdFoPrGhQqOrx0rbOlxutg5PVr8dyhR8wwcZqnKHjjKH0
UFvrq0wtUYtkIKTFs7Z6bcacW9MoeG8pMLDdK1PEKVA25C6GcRuHUuC8Y8JYOj1fhE0iTYKykaJp
KjJ7hNZ6DkbBynffqgs/o2IzpjD7a33YRtQQkTU+DrmS1IxxWca4szYoUxOOv/rFmsTOlDgfd0G9
ji75l43ZVfRbje8eE/m0m3SSPZdsBBTzGkOrRJE1om+z10tNSFmk0l6d+OclbJD4jU5cZ2V9Fvg6
mbQ8JEpUp+iut4xuSLATpnHYhcblr/G8mxDNbT+rC6RdXAhckDFgvWpYUoeYkuKBYwqd2/qs1a3k
0+m/i041EdLhUBKUUApKWlaqAw9OJnQzZa2HbwaPo/rEeq4f/jS0Weh9p6jd9Vqn2t2/Eg4XnAY5
xiMLwHvSPgtZEUMibLzvFjpn87sFC7qlxplwY5DEWQjPNCZZeCRk+ttiIN3DY15t3EqdOk01zerF
7mar4C4s4dJ8+4PpySbkkkvjRiaOU4Nx+FV97aNfHusax2dokZPOr0K5AnHcqdw5ef2AOGckDgVA
NLUS+dmsRez5nqYO7i6O1+8zsVf61itF86iNVMZzx67H+xYrIGgLaacLmxkHWNvwCos9BQVmHZyY
PDKEAvCIB8nPJiNIzKTYXJEv7GV27p36vNY8YU8iLqLM2JgI8iu90BVK7PNZC/RmitKp5IuR2INY
J5rkuWpMukYAuMp86+o4Hgq72I7PZVVyQNaXg4KH53C147w0/cREn9Oo6T2XhVt8AI6GxE8EUNgq
WbeNl8L4l5Y43ad4YXA5khQ57IjW1JH5nh85EAIvNRRU1zdDctQiKZy3GKTe0RzghjCJfSOM/3MK
sX3Z92etyGTCcg21Pd1PWbW3O22DhakfBNIdV1v7BvevSJdkb9UHiqZWuASUxVE/uN8m/ebuhnae
jYny/cIud4xfll7rFvWbuJWWVi/NSV/QZOUC0SXJR9kHRpZ7hATunVi1t1RG443xWvqeANFW6a5e
DgK4t91NSkRZqYsU+2qxU2nmGwJaKJaeejjzvoKSOgVEfYDsVXaSXYamLx+8NWvcSIUvcqMo4ekX
+0FJuzyXoh5UWf7yETeY1zQkm97TN7lwtWQ4Zub/7adzPl4BvXMVK/X33ydWbvZPsUpQt//RQMD3
PdM9KSJYRUxG6eXueMcU7SbAm8eTpIMLqsJsdhJktI9GX0Psx1WrzpK0vsUQwOLTPCJFXxeld4of
XAUXMl9Fw7ZfxCRKYNiHqmB/kIT2rwT+KjvQ47kLvUlM/JTVGrf6e3LIX7Gk9OWpb01NhAAPnrGl
bZKUkuL1SLzCN3+oCUjB3lcr2yoQhcDEpZBBeQHyxY990tTq2dn7r41QjQxS7+V7M1CSHEbNdaDx
REY2cpBfCaYUsbbgEQmcLGFVnGF+gOgUcO4P9wb9MuhIotnLqmdN8MBmqkfniHZZEGwCbmHTVOV6
w30JQp5d1kW7/PLCFqA6/Ul2YAYqwOTOwZZPZZv3wCRhn6kMnqdRgJyR5onxnd7+CeisSR0V1u6J
0RXXt/VlgoLJZwguh3azXvQp+bU9apJcBLFHvnM0L2NHG/yBdnYclsjukjQl2yPdyndkBtR/LBuJ
UZAa+uVEGZPtYmGR6u6L82zHDb8FCGNiWvfTQtQF+bp3vPr8JR4Y9+pBHbtAPcCJGTuHIlR8DWXY
up9/CjIV/BohYAcAjPtp4hpQ7lAkwqUiyI+ZeC40KUOdbgK+LJNDQx6+8hWLKVWbaySAUWlrZ+kE
jRPFjMozuhu0MXt5djl6HZpS2PU1VA84EZwUOSpO9NnwbSFI2B6mvMbbnsQ2jZBjpCEX6DpTgwNd
bq5goc+h8UjuRmE7+IYVBQCc/Qr4PIXY3vVG+V/mqR9noGHYjvYeBevMg7vxsOWHUFAtcH6m6jf/
ief2NyqXbOAmHl1UghwhRIdXJ15bBQ3O06ODAjYvEA016DgRkb3XHNdcvoTOyEDLowIOx5Ulqviw
aTqn1VcPDX7UCifQiHLAXsXNkckmul0EM6Ob6nOqFrJSq71Itw17FjZw6LC0/L1zAfHyLAT42tq0
9t9lnOJxTQlx+pF9KxYAoo35VmKu1X3lgYjcego4KYhm0LQ7hGpUzVmCUuzSEdNR7FTeWD7j15xT
vNRQ+OZbIE4xvykePcvwomfoUizWwC5Sup07tRBCr2gXmbuAf2wt/UfrUsrxBYIwx62zLZpvnCqw
QeBE1hO0EuNipjJsV9M6mn+wtHLU2AByU1iiied48thF2YPgfynQNOqd6nx4epXTHdL09zUxuIKW
yh+vhxEhy0pyMZwz5UfTkHIgkPlmzReEm/T2ekXdz306LZ56IiMja3T+9cMv3xH9ldao4yyIsea9
CVLzkB0fnICurKf7k4oIStmJQHR6lsF42mD5ImWECRNIVuzIRNrJ2DpKZHE5jWhcG2WvXJiFiXpU
fop5alu22rp6QbEwN7ApRokNbnqe8JdIJJKp9H6loxv/AIseKzU2fL/Pftzykp0vhoVXAyqwVNGA
7RjmjhsVXtxtaYwRLLy6bO4GRdldfVzF6klcnO/8uTl9exVy+PaWxIF8tJzcP/60scKsLP3SFOvf
xDAuj/rsD2LN/wUwC+xI2cb9zx2ZJtokFlPx1sSNyOYhBMzcpzupF/0gprAkNGW8O+n5ulDTPW2X
LTHQxesLxa22bqdoHE8UXOQ5Z80MITPn3qLz/w==
`pragma protect end_protected
