// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:25:49 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LBsIkx/6QyLjpEgxGVI3d9MHiGC6gB5CuotxSF6TuiK2VUaWLY04BtfRLqcN6hAq
Zbq5QFFFD0vsq8QqHVkvc8tazyO3wUexjHAOKfqamfy3TzkOaOwVF8OBdqAHL4hU
hGuzBdt/7WdFdMI6NwTY5+aKY+S6YiDsmDwvfrRRZg0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 36128)
DrV9e2AiWd36kyA0Hhk7RWLBUu9yBY/NBeD+oz0FhhTx/UmUr3KpTvRGYl3ADuGL
2f6HLZCQRht3LFfVsYNUQsIoKoKowr/Tu/Gt9Q+W9MsWPp+6/dnpMS8Dyxg0qxhm
Ik8QE9JGylOaqVE+mvdPda6yVFlbxhwK9DGk37iLxGJgjXGhlAvyuccqSi5CaKYn
8JMqwagMdeqPdLo9d31NjnFhjWXII70InGZxdmcuGzmBAZ2c5w0829+tcdUlp0zb
GhjWIUpWwUNE3aa6v/1PpmvLM7OO1ysELTvMVmbV/CGRuas35r0USO0BX61pTiNY
a2UrS5B54tv136eHBRWcgdyzDZ/ZkoGVscqGJmS4SXoGtXLw60LnkoFd9Kro2K7U
l7T5bilM3w1Z7YHLWqM2A7LL5+f0ZO5SgI6YYO506Rwj6O0GW2bRYrnmpB+XbJaJ
Vl8SYVP6uwDYOHVp481XlWyWw0SC7Lv2voonmLc5buwM2jJ6xNal+qR7EokuMkt8
Yzmx3pFJtYoAE0f41jOwjXJrTL0GUVzwc6PrPI7r8O1e5e5evlC787Nx5MwZGNm7
gLTCsbKiMmPTLWClxXTODr0lwzyHdK3bMvm2yR4YGG5QbOWrNX3GTV0/PZoTCoiE
B8+7FmV4kNr2tuLPFhUP/5FRnNsQ19zRzic2/US/Xp3FkwN6y9Yi505lUG+Lwmoc
wOmHUS2BLEKNtuWcKYHmG0UC4TYZ++3/V2wUbr3EBEpdVbzSbsJCnvQsQuu4TRmp
CWGxTYXuu8zNaRYqtqsG51BI4vPSRVVAuA0/yrwHLGLR9wCcFVtXOS8vfjNF94z5
JkZ4MjC/EbWjRSGJBI3PQ5MsJernvKpRxw06ydtOliA8Pcv0euqyQFWczh4QBFgK
uqGM80qNCRzhHHbMXSTpUwH1uBcETsYFyYVPDbafwrcIAiGxgWjyNJdy81nlrUNy
iUSmjqLg1z+XmF0dLe2IP0dA4+rCSgJyF4+YP7oyDAOtEQ5myYftNUe2Ml8U7vCf
G0+t+14B0AjbqVzB8nt8wtDD4P0KTJ6mXMlOOOScGbQNFCxLZqoEI2xYkuhVar/g
XHDhPXrsZ3pusU4KY0P88Wp3lwXb4Vv+RhhOd6Dhch6wAwUMn9QgS+W9077V+8Gd
CW+qdiML0jgKMmaAXrjEcoJOS9uhyWmOibGWwCeURwdNg1hiTpthugQRD9RnOeLS
oFWRf21jtS0eOv62lrPiT+F6ZfxrWBJAgctuImwWmZ4HmCQxqhIfeBCD2R1se8rI
6h8Ou6jWF5RbDhWwQVVB7RjX4oa2b9JkvkuqRxGWONexxc+cmS0O3zssDCuORvr0
iid5LuGJQeBFQOABV2z5CKIlT46gCgSYjPwhaCxO7H583R9oYwXVz5owSyWEPZ+p
6aGKhjbFQqPK7erc2Bo0f4xVBg07AFHoRpqLEmaMYN9BG9O1DvUT45YbWgDKS0ud
co/959bjpNq8lQUCjpVkH5XocSVhsDdfXKauDZc2EPHjS9agSzs9+S5CadwNqCc8
U7EouKJ1yG2aDtncnJ732dPENYEkAy2IlrgX0eu7nvrbHK6vgBpPTOBDXLvNGmoW
4ukeiOrB6qCTGzDgfQUoBlTFLdWMpSSeQveRuZuIyeWMlJhuTNqQv/sU9bjZJd4b
uD42R4fuHkx4vvaMHTQ/IoT4eAq9Fm1JNW4zViE1UaGCpd6XOLHae4T4pPjJ+O3q
nrn3GB0PQQpIVN3oPOqjWAbsOmcQHEkapX8yYEbQnK4Xk8Tl5qDHMLzKzJttmEYs
eqQbPw/zQUvS/FNCYYYVM0BzvVWVFWuAGdQTKGph7dvXLhBqnaxtrF8FG4TzUy/F
fqxvGiOxxYAsFrEhWs/Ti9xeHapd3N2ppdlE2cmBpM6LGl3mAi8sXu6K+fALq2Ah
8E5l18tb6OKreXa88ygYzOFe09dqcMtcw9oh89V95Cp7Mv8mzAk+gCOQn/at7AOg
d+6NZ5xctLULM/ZnFiii+azJM0DCV8jtnxEmcdkZFDZAuURzQIWWYTU6bRjXUMg+
j6RWijE4tDzP1Lsk0Rp71BOcmYHGKij2ASLFbbwTQ/4gVIFbDbnMjaI+QdvFF0Uv
J7A544e1qfBy4zNQThdVaafUByRLZ27UdDxro1jk6Wxlg0+/nxznmBsIsvMOFWdn
Bt812vZad645hTNj7sZEGY+l5gOv1EIbqIimjf9CNDm6DZ6nmulIG7gLvjR7UMpK
h5u2AG1otS1VL3Em+ICEl672h+sp31RDu43Ej/x7dQRPDlJt9FpjDrjKsjn+T/8V
qOXklrmVoXWkNBjFsfIQn6svzrl9FcH4SAGwkBqenijTyzotz7IdPR63XRluapDr
VsXkZHwGoUoOt/aTJpILxAaBSx6ApCjIGGFsGCIEbh8kJI5GcI1PyGBqxX7HFZJ5
PZr3kehkknznnWwTp60mtO6w57j2Wguj18w323hIBUAbvOHi4xfZXfwERmuE5PNq
ur9/BIUMpeiLxldg5zgdjRGIYJPwuWE7yHnlZ5pOzTu9kg0vD87tQf7zbYQXC/uV
xSmSYBvt621c0qgYLrJoasOr8EbggNekp4+ei7ue+z0mr9rOGOB8U51yuQYduduE
GvbMz+pwHDuz/fMz6dwm45fis5UR6qtyDvLRyJjG+27fgEgBXPmyTyXYGZtDznQ5
KMQJ96o04TodXRsy7vAx6G9NOToWDDdudVmETjYLaxBjEtFEt47ZDpZ1z9QsHzkZ
7wm35L3+7ibFiDUSOfB2i2kTmiRURhiDoxhDCB6cWREvPMw0P3qgDVmQ0P6KB4wN
fMRPecrFUjht+ITN7mW6uPm1e6CtCcDF3VeHjMKKzQ/ByqMxUbW/0+t7SDploTjl
R1tBGZK0zlfPXRRBIaLICf3O9b5fiZ8pC5YISXrpCCxCi18xBW+IUJ0ZOSKybX/i
gnmuxCrXTKed9MfTFOHPFzqFPQN/fzXBhG6MaTRqgOwCxY+6XjNwMXDcMwSDmdy5
HVyebIwHMHGK1+GdU6YvkSo3EvtFieAjbul7cswSBSLSSNTm67gFO3ahZhjJLOSw
9DPknt36ezNtVzmK/FaTYSoj3wX0n/obNTS1qo5pG7TyJiMrrV7m3SVDTmkthtIJ
VxFXD8vz387ckB8J4YVMEJSrLtZrP/3E2GyMIidglHRtqVGmaXLGZ1qDak6M3cuE
Xc/2CT5lxw1thHd7YrZJJZsOT/yZRv5dopyHtdtpl906E7JYGLXdADLzGEktY1lo
81Bt9LsrO89f38Wp/JeJ/DJszK4379y78mMfu/T+hmgjmZX0dS1dYvQRZHqz/6wq
GQL7Yw0xLn7FZxgT9TlCqmziCgZl+YuKGlG8NcNLuF1rpxQckxzHXTcZ5RUqjzkl
Hz7SUmIjNe/79y6MmRO/ArgE2g+mjYgqqveDhGNqq7khDjchZ/nRZWKTeaUmCp8D
f7Z8Lg9cdwGIY2e+SJdG8hKHJ9TDQbEca2EZ27RBYB8pdR3wkTaIDJ/IaJM13SLT
xLqIL9JJNfJW7NKSd6kzc2Cj+ZN6/WbAPyU1nigUjxgcZRNwiMBDRrZaucvoOA8P
ueahbTtkj3ZWsvrfZv0olK2ZKY0KLQNvwZq/PRKXSwZ9nN15zDqnHoXyTA/S8GRg
n6E8Li1TA2dFehra95chydsucmMEuSZxgbUzYiO+K8q7Ui0JcemnuQ/n4VahB5Dw
2Isf5gJdGuWiWCwie3yzfwntSiwxq3+2ip5GiEPxkpG1uC+hf5/zkJYHgnvFdwOv
4GApmvIKbl1nQ37HRcoveeLIsVeknizNToFdfD4/eiLtvwICHp6RL9GD61jn2zWz
H1sA9V7EDipE8lzX9GnWk3pKvYIVOj/nBM2eBLzMdfa7BWJgatrSc/61/RXoFb0X
EXBaDOj2LuvBL4DYdvgWuJItNO5e7vL0ItOFdB/dl9lie8JKT93pwo/Hm/5Fu3Uz
jnIrcMjipdAiIIV7XewtSeknctUXh0IJI6gIh5gtnziCBgJh7MmS73/VuM5gJm2U
sA3sv2fBSmvmjdTgykCP5k2QnJvn1/tP2U15klJ9buJ+cNm5WpRQUFSlNcxYpT+n
Q0MjR+jIO8xdJ9SSqLzJ63T9O2kVRs/PfAGJTZUxUg4w1Dd+1ZBkgohI+TB+f+KC
7LIhkCI/C0MPwDnlHuJbuGAY7gz3hMrrDRrZuWlGJ/N7C7aWBci3xlU/A3b4EeCv
8V9/FEeEhZEQMrzDOuidZ4bfEeHO+CeOkMImrbLQBkBZ7KZphFWiFTygHO85GzSF
rs63BWI94UAuoSYSOjktQUOotVtfLx6PRahBfWrD9GGaPgeu3dsrxePZ+5qNaUAM
sTvdPIts9TbjY869YpU0Oj/sI4hrFvIfRzkdfcn0nNMZJXGiEZKsUZQ+G+Bkm4a3
FmG3zFjHNErnUfWzY5eT12nU4CWsTd7J5WwrqpnSlA91VwgVHalfFU+H9keFuuVy
ZoeRwhU0/0XXLjDzoisCCAuTAoDV7XIX6d4PeSSKTklB2c2uyLa4AJpIOFILiHsl
k84KtnNd9D2zcU9kobvSl5czEB8L4Xy/1yap1avT8bA1ObpJv/xLutc5IG7m+aq1
CcQmi4wKaKwH2OruazaXcqlgdr4HEnmLfxmj3b1eRiSgxs/OiZfqfsbYiRTMzMBP
ZEjW+Y9pgqpegkH1/cZV1vOgQvxZBJq3yPz0iOGUAS6XT0pWHPEbvhnvhUU83EEx
hICbWEtXVWYEsjBdM0SOc65MZeswjafyon0JeLFiDm5OPY7CrNhHAScgigJKxBgC
CFhTfM0Sx/bFvvYOqqWcFI1AqUUMJ5wUGRr8J6+OsPaCSyG/Emqmq68qeEtjfmTT
ZjMnrUEj1aVq24UkxC56z2psKRF3y527R/PbgtqFxkpLk8sXNo9qsENzXFcu5/Tt
7eAuP9N7h8iJ33/E8TJd/cvkycM/PXI0czfux6HCHgo4FgNKGnfHPRAMIg4+4ro6
BuEWPhyadxtDFoAlJEwj/HoB4bOgm1hrDXyVzDB2YUDwWxhWsoffybWRM5TQcwbO
385iJec8czkvdhgewIzHa+7VjoDmXfzU+2QaiAhIN2+kl3alQRHt66L4DqnuJ4QX
h7TrHjMOUaZzViztuZRn0Hnxz/aZxjkIXFho4eDO4pEFiDb+J4e+yd22KMEbLc7R
V6mCb/jjPO4sShm9F+VADM1BPHdfVUT3cUe2h/XRlYy0LNMgllkIvJx6EXPVQrf2
XrlyLdRPSS74uhsDniu4dHOHH7wiKjlukc8H7GOQQtJJ9H69ygW8pja7qPV6mcMo
DZ9SFRKF0oTRTWbdBHcXdh8sY+bTs1CXQqOy/OWEF74GTaLYoc0txqLs9PWR9ckq
r7j825IVBn9F4onDxSrMLdi8JFkimIZWQDS0A+GnsU+fh2MVx65LTUKlLlvkrRT4
WxToolNierXN5YP8B8Ehe1V7hUn9eHxxuABxjOi2+zCwKaeN2OaD0VGDyFBD1xLy
rLmj/J8+F3/wf7sMuhsAS0qsFP0WL5ZQaVuVNiYO1lVaGpjDg1SZhC4LnJWUijWx
yntTeib8n1umwiaBY1g9yL57pHgZzerwe3XspHhyMyGfGY2AczEPHJpgoqXko1K9
hftAzzF7vIziWBV6W0g/7WhyTMRm08hk7sAjN+cFHyN4YTymmnAx4mdHRyHvfonB
CrNICnHXLo81/9ZfkdM+7JfuXlDMZSvhd2fwpS6CTWk0dNATT2MmT2ggpbY4cnTI
RIHJ4ISjKCSmsKF9RF+Qowcq7JWwpS8dAnBi7MoJmIhSqSTd35fdZ4vZM9Su4flm
qhVQakrbGu6Ee0gxfZN0q+GNwmcs+A6KJzWUjhof4UI513yJ6kX+YjT4LAzAMNpd
yU2O3cy9j2MGTD2uCWdAk4J3vrZOruJNek1bTZOGbTuYblFMolq4OKrG/S3/RKmn
h9FRhhTZC3DOQGBvXhVQa3KCAOuvPDhoN8EOk8tQ7QkMhERbHYSPvP4bTu5QOMp9
oS//uXaRRsYr70QxTqb1X6U7ysCjhWF58qVV8OGndhY5Iq74zq4wZ7RjA/BRGEPX
/s4cWEOixO3sRHbeIbMCLQkQmqL5iA3a3tB/fOxQ7OJP95DUod3gMtSiUCi8BQqa
ogFqexgDCOmjKqSVEQzbzrUwibuslXTlr2BoHEO0Jr8Rs/plRLTaUxWzq9hjM5De
tXTbEqYzQMsTRccgkpL3pg89+Az8BtD1dzTVlm7O6bgikw6+p0WRtfxlKVUr/25E
PmMAJi3HkHj/BYPSAJ2IdNZfodEGNreMyoHNUg48H+26iH93FzCdH5Cc+AVf7Kp8
vhk+jW+7gJeSQocutoG9sprmjzxsSwBzTZdiWh+Z8QokA3hncn74gQUhdXa0pa9X
64uB/D2iC3elWbmD8JUCrZukAbnHw97ZCNFvfJIEfssFo2nY8X7uxhMfO5ZhXWPY
Cb3zNSPJ4ivZK3HhhWZeyM1uohrY2CHnERSFYU9Nd7teLtcLylNG6Hu2eDMDcQUJ
+NVQPXn32SK6J5pae5XyplS07mhOVI+aCGt10psDnwTRASjUlrfis/VAzO4N6dDX
NXhx55aku4pjfdejytzlUHc3D2lCWRLhV26J9mzJuigAJV97U57cBouFahOC88NQ
cnIKgyMokyzlY2IcnjTXkvyKk0jWAdhJr7yGQ9dguqF1iDg9pwZ+yVLr4W1qK5N2
S5wXNsZ7P2awsyVNtV59bLACH5sik4XbIdj4nDm77sgJKz/ow8VsQiMGoxkGU0iR
YTOMddL/Iv/aNbD4OBk2dlYdNfC21ssZzGL+hp05InvZRmfEmgSYgaSP7YqmP+aC
J3iV9jgMv4uzfSPR9b+17ydF+7Gdek2+u+lPEes5TfQvRSgB+XFsXReSdypnBJcy
6C32ZAOv1odavUPTSTHPQ55HqPquUgrH186LiGWLUvpR3V/3CA7CrA/A/DmcoF5x
23WYoqQuxKwafZcf/sSp1uQExO+Ex3l98kuZ5hXgZLJmWENYwbK61PGH2Gd1GNQz
fE/ho+aAqkPe/FIeXOLnTb8x0GWyAf+V0f+HflESeQ5/Xr7ax4fRPMOGHwWBVvS8
MkpQb9HjnezZVOZRbdovYomb6w9wbJOahfw3bdPr9cLsAZNRRbrJ8Cd20HEHFPTJ
bkm9ZLZ/eFmdTVUTpF4F/4oX+f7GUGwVP0S1Ju+f2sVhTvZ2xxedcPeyQbOfm/rR
gQc5D+cfJco9Z/jKvpR9dn9qnB81gbSym9MAUyy6JUQqPWPGPi+/fLvpnsF2GDRU
D5taacfYxRHtADP4iymazI6TAfj9RdsiFsTuu4LIVg5OzHophN7yLlo+851AHjJI
TGp2zYZKDDXivcET7MZv+a19WaRbCE82QR7C4J1KflwaBN33/fxvTjdprMFariZs
USyuG9uycTQWpnaLk+j6gH3koruLds/T+G7kiMnMscRiqrVC66mwsplM0h75XYcq
zhsfUkpssbqjtY8lHxnvKPDTSeeHm/loe0gn3XQFskehwAb0UGTa2R3kj/EsWQkO
wvENqUuAmXk2fB4/1ojClzbY86PWaNQ8qMRAwjkbb7PbStUDu/FCt5FeVuA1M5zW
fapeazQaE0N5NOCjfqxJ94C8rpfxnv+EkdK0Z/iWWOiSBp3u7jmCxJNlFssUZBOz
saYnM7Ug3Hl2L7M6AYWThpzK5P2g/v3RfEgMZq670rBdZ1oQOmsMtpWBxKzmGhp4
bW3HAFBHvJi+cqCM/TmhSg2Ql7ix/3qnrZa0izMdMhNBcwNwj30N1iNPuHmdzjVh
Gs+gJMpRDgiOkqHO5cCfGBE+wKEt8MPtMBA9dkca65+HolCTB4jr9+w5JejNGxmk
d3CQSpNlyZ4gr/gaAcMLoae8ARYkdXuzslntB5VCN+R2n0h9kwy+sehOCdHEGRDG
6HB/J+Ek2k2Rk2ku4iimjfPndi2Z6S7+xtdpFXjfkmhBj1ST06S2Cwkk5yZ2mDqo
4siXPNl3URNMEzE6FYh31cPKKrbossrtKUy8m6Z1exdVKw5hCRWSBlrb/48BMtfw
vg9dQSlT/TgWq//604+l1EWyprVoV/ebyc/kyjHjDTqkzp4Wz+vTM4cyoNeSx+sq
0Hj8HzTABFMCBPuyJ776h4zMLbAauIH6iHTJc42nxLtncuKH4NHIamTw0EGk0x+Y
xqEaljjJ0pYQ9fWTUlRXExAPYF5tbAzZqr6JqJCtmFdtN2nOaSVFeKABKn2nrygZ
/XmDr5r2LJs5F+SL/Zz1h0chIP60Oox9Z1j3pYGvIevu4+o0mUDCLCGN8+jVl7Ci
IGJfRSECq/hjyFHjfrEEd2DkgxJiCM6h5d5O7vQjUdCLbZy9ByUih5eotUtRveun
ltct1CWqrmpyKzA7SFqdqI/OIr5NP4BIvNwbFj0qvNGBFB74exwZpjBIkGiUgDwd
ibK5jpQfhNaEnomzHfULpvLxnTzyCEAeGuNNdOq0wwGydbRXv77ADNkUYjNGvF6G
mcFQhKxeD8Yra3C2r7ebF/XBn1+o+EleyOzhfW4X6ihgHfobu/uNQDZuTp0O76jv
gll6EVR9U8X5M9xudXlTrXDXcEQv9syIej4UpOH0W1fZ7ZnckeKa6iL5iraJ0ceY
nRsP3xtnIo0JlXtzGMA1dtwBkJu0/AlU4PBn2hWzfyf3/0ymu9f271y358aZQoub
7VJwvNrqe6Qiwg5WNmeFZIsZXsd1ZSgb9k9SpZM+BxfSlLXJTDKGAFf+8Vs+nm0m
iCKNeEYwxbSHcwSKPVjkPrmFf14N0dLP767DgJlcyGM1EJSkkgCgD4jlCycHKHd0
szfEdoS3aMAT6Z1C+omtGqxg9vC0BEF4Pvm5eOP/b1qBT6Kj3M9lQCnNMeUm2FJO
Jw0rDkCPXUDVaDNdQq7V9tugg0SMespGWMPNmW3uDDohzCSWfYGnqrs9xiZNVr2g
aRbMmK0w1zWw/eoogkLqogFvBSYJXuAIe7TcJTcG1IAwb33NnirqS2qeBN7QtMol
fHbcbkUywM995FJnSNeh2jP05AONB+drs6RTXO5GGhXwnshdsyyawGYFhNM1u1OC
E1EuZT5N/d5gHvCDLe7zT9rSOvXovWJyBp0+SJ6M0yomUjHYoUBm5zbEoBcmfRfR
6Xtyahr/ZEDAq6YJ8ixscYNKkSqCdhld7NWlaQDl2s0Zp4R/zmVGNA/bc+gxlENC
rVjb9Svs5Z/dfMYSiPFThvFJabZIFc02930BuMz6kChHLVPsHu3sCSQ96pitzPAq
+FP4gkdy9U6X94AqrWtt8zhezyj50G4pdyz/WL6IGyUsZ3GoYPtpmY9l3u7b7MJx
hGDSijEk/0rXFMtggSD2QAN38uykpQ/yATlpTWyjdW6nhKzI8QH/2a/U6VB9Vcnh
8dOM8byRThr5JxpMVW4eQxoJfQXpG0d5BtmBDfZ7d4DvI0GNcHq2MnwclaNMA6Vd
xop7SOCuGuiBQHw/pwj+1GmrZINmILcPDICTODvHLzJTkLhkgYIAbeRa5QZmVdTx
/bhz9ahPf1Ong5RZ41cAy/b3EsaXSOh1axM079aTQw+7VZrJZPNds7t/8vwEKpBN
R44tj1+EMjCuunBlz2s8lCWXQr1ZGf+BFQH+crCN9Ku1OoGs1hMnVBffC7h5O5xX
ao7UPOddvqNA6KubA9kr3pVoxyJ9BMw3Ft4vZKQwH9Xbw8ziMzoEgyncp/Hw1hTZ
1b0LfG/HnSlQi2Y6ZZN5P7UHCIhrlnbNdrRKqaYb9GN6s5UdIbihIWoA1EFn0HjI
uMxFGGLSbag5DqGCvcJUCM9KEEXMjPw/LNNCFcPAnRgqMmIe2Cg3YhkWNBfd/AQt
t2x1Q96NDSqVRGnT0JvxhELUnQ9eOoESJlJ1ze4mewg7/fODDLS9wte7iPr05CUs
HJc+B3aoPCurBZnxrlBAlaNicVGLJi2ewPAMgZkDyhFmEHTAvP3+lu4W0FA7pylq
KCPgTm0WKaKgJbljWI6hTlqc+bIc8v8dGscosxnsGVftkfUuLwLaV0tCmiDTwc70
b8xwkNZT4qQgxRyTOKcku0WIf/f+/k+fdz7oiuXS4XQmnTsmwYaOsyBHDJ961lx8
AuE6/UPg9M9LZcUQSdPKJaCUnwG40zJvHBO7V6wZ956ZhwqlWKKFQU0anWsG49XK
0lOjFbiPd4rV49pub1QoAgn+4ilxh+wvupKETUdq8BQjUMUrjAR7SU5qitkbo+KX
ho1HeIwqKp6hk5vx8nF66oK0t/JAg6duY5DI1nhxsLL78UDY0Om+v89hLSTwB9+0
ONUTtpciuX2GhliR9YESq66qSzccfA2A1CtRwlkdwkg0bXIUyVrq4iIY8ilGS7Be
RcLy/5tg1Iior1sEF0wgUNakLpMWqR4b+FzqxlCktYRe0NyWzcvbZgWyHUGROvxG
Wp40nShz24eq26k04DkbAjDIx/0nvDC3SIxk2GVbNNm5/dQxEwVvxgMIGYn93I8Y
sSCkA9vyzS32/xYdv1/PxFZKyP3AKePu4gMXb+9i7ug4ONkKBCw8Eqix3/5MADos
D0hQMwqwWTWqFhiih/nezuZqEDvQZfBWSETrbbCvEe1/nSxxc7gpyQh2bg7IEuyG
jeAxKKEGTDvP8+tGoGSH75Lr/4Weo4rGlLIGneGDxKmFXUSlVzYIjGz8DEPXdv0/
UCax9PNcOw+6QEB2gwNbsgWmomrnwU2fyGjuwPE7Pg0j+OxeB37ybyTKwESgGv/Y
2GbhPhzqUt5p594sY5k/F8P9qQsbWm34x6oTHwLmYpKXh3o85EsMXr66NJ3NshBO
F4nsOqAF1QsV82rJhqedu9xQYWsskShobMXiGbXal6ogUIINDWgXjyBdYdw3+psv
ZTPn5/o0NoUhzMLEMP3kniPl88DgKfhULvAUyLgMqb3+WeYKCYk1hZEzjxOfKehx
gFeKcGLwfkJb8kubwXYeRtIGX2FDuq2N7jIJRot7Z5Na6TujL8Jvs/gjRqzNPaYp
N5nL2gnhndl9y2pFV+1QKEobLFq1SWEiHxLijrmEaWwO31rgwh8UhSR+/xxFhBEl
84RvzRFboz7JQw9sA9skCCxQWk0rPTTSppCcyROZg6Y73Ef4kp1T+8b2VhTUdOYu
1eGtr0HxdeNfSbXlqobc7QzE1h3jWnpCD9C+uiBVoyPGuHuixHAG7BTf82NES8gu
5W7jVTkaC9OWQ+m5/Nzv4JaR9QezK9qPYy9f+/3ZTQ2ghaFf/g4vaj2irUr0Nn1g
nHHflNyGUnPVTQXpRAfQRNtiI81TTl7DHLypWpNbwqCuWLRM5zqZTJ7EzoaK+nsv
30KAj/xyBN+CZq4KKFQyBhaoZ2aD1uo9TnA+5mUx6gGQeOEim1jDyzwFXTv4TUSy
9msZe4cl6ilk+Bz9W2uC+ZDedo1vB9WGNrt99WnCNaSjUHsGOelsSsiBXIf9/a0+
lSJO6JqO9O/asmIp6On9pC5Cz7ZqEhzbUltwQ1TBvmAXdbFCu7PFQMc2i4wblI+A
blniw6HYYGYmiqTaczWvB6BGhJpZWmdbTcdst9k9gUZU8kaAdqVSmH+WsYjgwSIv
6j1HShT0yNQW773xaethS4q4+YkyXLQEeQH1vTgLhGByDs64jC58Xg5O7kfT7u8J
ouS8oiuSZKDx5S6M/RKIgxgjNZUg5dDb3Kz3uRXdpA+OptDQlIcz2vy9bbVUICto
lAaEE3ls/xrObBb/27UIMrJHPJHyKzt3YOVtMak5sbOGU2iPkPoRUxsbmnkBDoF3
oSfK61SWBii463arvXfFVMGZWdMLQKAKa+X5bC5tP1wFWUTnDr6bugwQajQi9cxN
cEm9Z2RdzsPvMGBdx9nz7laXdRy9ik5aPzAm5rfo7s6hA9cplfQaiZjdykRaf25G
NdDVCk6mPtaZgKtq16287at84Ugg3ZK+ypOOPs2yIwRflKu+mJVGFHFSmyPvumk4
TV7OzM5/YhCFKcfPjvASuoHAr8psUotWuvdl/tu4IBJNFEBD+cNqo9yeMQNpYYEJ
W6snhCgdIlZ19aGI/V/anZ9P310hG2uxgD+gg++4XkKOJyIUQT0EX+AZO9IXKPjK
rHuOO8zWzASI6R+O2Fwe/P/wzbfTVvUgYJgcz3kmO51li5dEfj+FE0JkwZC7Whd7
M0A0iVavnOlrNoDLWGxEYmpYUXpv9YkUn+PSmbAIiMbgscnUKUNf5tRAZ74MOLc2
IzjB/Z7TnHVGteqk9tqRpWLLK//eJo3qT9S+w6Kas80PrCWf5gTxTX8UltqJwztT
e7xTwHcJdyU6z5kXAXt5glnbZXHMQzg8LY/GP7Z0TmZ90N5vevpMVxeElqjFzkzP
DO8NxrCSUWmy7QKo19n7EBuuqFoJ3VNgOwzwLdDk0MrNq1IPuW9NMrpnFBtefxxl
zE6cU/ACv2m5ZW3mPbQbOrjmI0aXYZpdCIuC9r7WaBYhzOVC7/LTb74EnNmKkxwE
CS1AGF3KcJnvHyozSHvJW50uo8dM8kRUGULyyX14bhPl2L6wgxp5XgtViCDi9xJZ
1RTGfZRwZkg7259HXWBPZIawRcC+c1YxgpBx9YaSf8O+pdzra72+KF8VPLkkOuE9
2Qujvdq+1kP5z55ggJKrC5KXxtmSHyUKWk3LH4qSDmEBDHnR1ObE2Fzt0jH/fdqO
SumclncPyNPj/Gqebw1yq356eW0GAsim++ORCifz8haWoH6N77tV8EuvuCV1XkTy
0p2PNZFiB2h2arRWfvMLmHWtFQ5St7kQjB9LDSzcmXGoSd9NgcS8gIp23jlF/Ogg
gsA3IUAC8razNlR8YILiUCI34NJZ054WHN8DHrB/ze92KX7C0uG3WoGUQjUmik1H
DwxWmRY8MHgSn4Nawqx5+AlLLMqIwGEXAQaR86laBESo8En0Mkp15OEGXJ9IeGKf
CcTecVbkhQY4MTwyQTVEu1L1bL9k6XMTdTFcAECSOBLaTADnj0CSecA8v5vcd8YQ
Sp5+MeLr6/F5E9kelSAAaalP5E3m7HK6jHsivqXjnQMw4MuRf1QEphVOI71T8Srx
PnPR+7px2uEurFpPJ6Nqo9jaHDv1Vyuo1rau4PP+o2XUqYAD8UhFTn1G72ZxXdyl
mfIMbLa7gRHN5DaO5F1nwj96g9yhkLGIi1inAr8yxvQIBWz1HLdWCM3/4RTvmGrk
zrmvJlpyhgyjY/39E+s1qHWODwaaow7aQURpSS3s8keuLOiD07twRqGl4wQWMlTd
BtqMi0/mgpYO12m/pyZgXMwjy/hItYPKCTGHNQ6fu5OsAZ+u91T3YeJhXW7Sdqo9
M7rzaBhxfpHUND+D2WJyNFvoKFOt2uN7rA+fFF2pFAd5Elt1siIRhtqwQ9keHsY9
zZ1MAbi4A5WB8iujbhLe/Ctc8Xytrz3vK8yeOfM81okXq7UQMqba4cziwKLjXQSR
UAKRaZqj+KPlAvwQWKMAZaCUkKCyOzjptp7FdVUu8JfkJy+mL0MRBqiCaQQ2/Uan
Jv4tZlMIxYCFcHP+puTPfS8aczJUqOGl/yyezX5l5MSIYw9i/abuOabjDgiNT9s+
VW6UtKcTzaVMeJ6Lm1jiMlEDUFlmP5haizzxKgEtPP2fnyqXmcoJAVlArW6QG4lv
TB9a5zP37pEYeCiTiz9SGps7nM6oQNljerdD//w/9ivvHXBLAMqFwi3BNX2oa3Ad
sIFjyHASmZZhlVsaLq0VeC0zpsVZRr1ZcKMD55zxaTodL7bf9UTXP1bnUVdtSF2z
THDUuJP78j24ZJDld88+oaaHlOxOOpbWpKe8j5TdF48XWzGUbWZlSLGDtf+EObvA
1zzle3sD1u0kBnZis/4NetTXadKEZWHJ/S8Usw/hjnQp6mccNwe5pDoIzvQqYkJq
vkM5zf1I7XxfFtt/VQ6CXVPWbnj4PHud934dTkq5FEAMv+wySb/ED/iix8929mh5
NXrfl8Wmhdh32nrerjA9LtUsM3yMI4xrswcL6OS38fd2kkL8GV/NT9kjgKt1guMk
eWVMZq2PmzNHExcd8QYul81Zk08qOrBDvwEfKVDU129wGZ1yJwjs0qMsuSOh90hn
OqclwT2xvV+Kq77F4pnV5q5FiIkcTS1Qu6aSURXI5aN7Vr6DkjczkeS7yCG7pqQk
+eW10+nHHApSfV3ChWQljjphjDF9Ou+3GjEdyZnZ6KC1k0TFNdU3Pt7XaQiD05Wx
VV15SmXaQ2owbUFi4clheW0KQuVzrQybvEDejEYPhHS81lvBSpq859kmrB2JX0Tb
VQzUX/xUmcqzEq2TyD2s6tqkq7fWPdEUv/QqRzPZ01lJKDjOdWnLj7eOinaKymiF
50J/09RWpb9LvA+jWZE4fXqYv+222mdFRvaQOfPaDxykTF63C+z594neagukfJJE
62geDEQ8lnow+GfZwoXCB7mPGj5g5mRAOLyvDK25PySUym+MYdwU1BYXDcS1FDye
KTVOEsEbESnxOXh3FW0IlSB7FTp2pRUmlRYF3qk6UeoIaGUO5lhbKFaXtmWT83Rb
byQWCmj2oZ53LNY6T1hYUTYdhKEOHFluLj7/Qo6kNfgJdSOxPSO0ziEuMp+NVjfU
FZF0ZAAE++h0lEtbcWp0rGLq76YJE85bOVSDuWxWlOhnn20oVNtBVs0tOR8WnFsG
CkJmlDjjqn4wHeBjord/P0DqCYy4XxcUgnBkGXHkxgNjtRV3pS+PxqCJZJA38Yxq
G/q5tiyXVuZiqT2Z/GzwvP+FNri061JxybDqLaj6whdeTw3VSrAfCuAlrrw2mhx0
sCXdM0FSZalpPacHjhIWY46HpOs3d1oceExFgX/h9256IJNLg5lxUdk56iVG5SPG
5UZhs8kuBcf8fwdhvLWLP5U2lZvClhKQ9kschMm04zSh1aid7EGWDIIvK1Yooxgu
OHmogRW5TQ7TnpSEGmffqYqcBWxaE8T8KXwP7S8lREOWNEd6NPKRFUj5sKNSckr3
tY1RMHAyZ8gX2lj0bJyzHHNEwYb3Fm4bIbqY7oZsbBz/8dEKY7JjZ7RA7s+i5knn
+jcCj/yeZAb4M22NDZvj5QQtBNpVAtgPEsz5uko1HyWKrw4HY7CDpnnzbIlaQzqY
6dFX+U25yo5FZmSiabtzqm+kPeL1dpBegwbwtwcflccfSLvZi2of62iCAOQcpXaU
UmfZIWwJP/TBnIViQ80qRVSm4R6uGE2kvgo54EUjlanVeJ3wWGXWRLifaEH4fFtB
dMKWL2tizIzW8Y+9LgNwc1byLiA6IeBSKVUlwlPqHI194kppttWtQiIA/9JYz45s
63PFVxK6J4/M44Qxnfyw3ddr1l/8wkRu9QgktIOhozPG0ingmiFAKIpDx2tEc1Zd
jt421LI1XhsJ1xESgYK6tGSyL6iBtIWjn85hJX9zhJYkW+/dcjrMPkY5V/WEDMjT
Lmsm5r3Z3E3f8qYnTe0OLrW66yvjxoigfRR9lma5s2Td2md9cIrz3GvKEuSzbI3l
toL8ULpWpoK/S5vTdpCQa2KYRVWKXu1MYGUvZFznBZrxaVgmGTdbb0oOTyfsphyG
njjaHj1oIfIlgwjqeCHYWf/IxujC5GxbgVtqXeIKYFWT4HSiaTTgh7r7h9PIGuF4
ZwuQE8tCBXY3O9QHUrx2b1IpoET+Up3kOQH2AGY3259LNmAVs7QjzlPnZZw0/Lna
H83gGBfNz4pgly2AjiZajKekghjzfuXjxvdWrl5AQG68xY5KclbfczNasBLBxuHM
4XGhwbzeBWIlucGmV1eXGLohkHZq0nH15U/FCc0BLzKaBC8TYzzKaPTcgeZAaf6a
DiWz6Hm8cMlvpnhWMk8OOyZX7EPJ7qimdtO35jezbHKBGGGmopcu/D2DaTis+KkV
LeAOFGMO15uIqhIAkQ0faSCZ9YARiuBZjXdQ7fOoPX79wxW6NcMOmJ2GH9sugWDE
+rGKMPXDApbnVpDT2SYLzRcLkw5J9Vo4gYXImZL6+F+mG6uPhtByTMTFB2yz4Nrq
p7ttohXUKCDq2TCnP+P31h3ew81Q24NR/vX/8lkVPSaouNRoT7AC2/ZxRnCSyNgH
vXGFuedrzJZiiEFH/N1yJAjJBoJS2Z3Z/BgT+R0hIxgRchWw7rMZz7bMOtg4ZwMm
zWAeJRiiyOPK16jC4EhDVhLv7cRARDsyRm5iWL+OCz4zEvjJo1+gk2/vgcGlKNjD
7nZArA8if0u5BFgdd8GYikKwteBup5MBbRKGMxE3qOcQ6I7ZDUwMQW63lsxatMr2
uDVlJIy9WZXxKGRkpm7YtR7yuSeOUo/cWPuzoQftYnienRziFtOHHCmDewu0pdQ4
zVvOxQEqjot+ZuQRy9+mOUJpr6KahYPK9y3gvWTT0NICLjPtnykn55njnMKjePPB
VhXEsyK+X3J7moJNv09yBvR7CJcyZCQJsGVnk5h9ROomFa6Pg3U+yvNmWvFrN6Kd
tytyZPCI7726y8iDZ7Tn3PJ81d0gxr7jw1rskpSYcqbrOIIP+WE7N4WgsdA1nOv4
a1BakjKTWUi0uB2gLi3V7FHosB7nABEVpfyCQEviInsaWl9mIHlFgSs/TV0BHTeQ
v1M7l25ddDuiQ9Ti64SdRp7SxelVl0jsb5RU10VGedFzk/5KKSvR0l1xP8DKZbmz
54D8I+Sk0vOD0M18MCAUbLvkwlxpPnC5afHFNu5G37mZCvXgXIrdm/8An3QSq/2s
a2/bcD12e9qHj1I06biypQ1kgvgEhDe6Fg4E/fnG6KQJnXg40q3TyqSU9RW+bb0y
mpq+2D17COY64kr49R9qCB+tfY4UvaaFKPYPQqNPdu9fxSPZ4ofP6Nm15/0sZWMy
jZ3cDR1H5wk6Q8UMkzhnIyXl05Ja7VOvXFd3AzBRhIhMRf4YRKzt34qGhURBByUQ
/45/I66i9GAUKRQPVtv5duuaF0c2824Dv3M/C29a/y+KD1MXL1h0GpfBJMWIvx2Z
mY5RcWu8i5wwNFPSVBrjFku6TBkPgEJ/2/L8yX2rHLmRtNYOUuIHFwE0cNGnCGZQ
9CA1+HeaTDIdkoh2eFQfc07G/2PlOLjUVyfkDoRNRkSEwyUjlEvOBePQdRJzL7wg
z5pGVT68nSwNOwTzqr+VJsxVdTc+xibedOvwyuMd67gO6yPCGr2p6f3Pj65sJ6MR
o5/np17sUkj91w+fjmoKqLLSuN5dmI8FFboueZ+pzvYbsnIEHpLKS1AgAiu4G/Ex
nv30fM4WIb+pkGR5CiU03A6pxKtDdh/SH/DOJe6+/INYTBe8fwZ0F1EDnot8BR8m
g2zDUcvyaqFtVW0h3FfFlemftIxiqVIbNhRczfJEuXopKvCgLlS8aMrzRQGSieHw
AoJIqou/OB0SK5QXREKZjpl9LHkEZOlBG7aGc1zdCdUNWRCUdHRlJGBNI81QinQo
+nnOMU+FSv7bwGBXdt9+BGGQZ9AJr51oW2DbEce2pR1u5cklRbn5rIYXtIcAmGZz
c3vb2liCYmXHmRKa/4fqzQ2lVVBtyUGfUuRDRFc6FVWui7VqNBXUEHDPao7IRfaT
eXcg2N6baaJakkCl9toUyWqPvKNinoApdFeF5tDsdhH9JdAJH6va/yKEh7DaY8jL
8T+M4XEzLJ0gz78ea2NIuRHEBKXzq7RwGmGq0sERSVd/Ao+SMWf+IWadRLdV6IIu
+Iytbg6zI2Q2fpDsF2c9cEaB91oimFUmMDkoY5MSw0De56iC5qnxrSHZCnM8Sc4k
UIgVaP2lWFiSSiMAKGWs7YrxJY5fU5tVm6lQC6aY+5PoyBbFpjTvHVq06cjPJE6Y
7V2e5dbR8gkxm4IgLljWULqioCZJNbqRL78Gv9bc1JFfPBMjK055ZyutxFx4DnJs
bzdlw+ncrEuuojPj8Zt9vr4TFid0VhA8aXIA+oQIeCyFS9hNMbiqNbGQsOofhkDN
rcPZJA+ia/LYH+V3hEdruoqjqTTlBIg9BrB+kxgyRo8IvJiRhMFTXOOjLgAso4CU
FcmCxOwBN7vM6AaJYZteVSZPEfueNi/XUeANG4tDznXw9/VkY3n9hCNMaYn7JY23
1vS9ABHLxYHht36zrwyrNnxVsw96+CoP8zfYeU+UMrSaWrjVPFpdTUrjazbxS8iB
U0LvaSQTT/m6ABN4PG/vLvF7TvEV31m0UXcfjH9KyjCoEbKYGDYFOkRgqXsLLicu
RfDxkHDPOjqUoFexJhAh0r4o6LbCV1HfhbtMjTeNLPuazz2nYDb17z457uf/oPWC
u+fWavE4lyKcUIab/XWPxefIc4OPa+PBfgiNy5hGgqV/gsjX/aAoNG5exNyMVkoc
/59NBfYNEHtgQe/gm+9cKEgLtMIM85C4Lvisji/duHetSYIL2X1f1zweAAV+ubTP
m+cVftP8/ucl8Zgo4V2t156jK0/mq3iNitrfP7t2z0rp2Y5+iDOz/82xA4/vTZr7
ZFBkiE6wgNcyG/QtyPg0YtEByeo7Si/hEg/UI9eICXWWGDrF2LbCrK16COcHdtwe
17I14xTzIiKd3G28f9hpTqWpG6qbgjmn+uHEVqt0aOLs+5RST97ZLUorUxOMf95F
c5DwKGUPi3o0PCfdgTYE/LaagVNb2BiBwwiFclMCiwTXYTUN8gbia7IVDnqitkec
lyzpFeG+VoO9TXFW/zD1Kdi4sMIXJddtvXWRbgJPkeacyqeAxNz/mPeAhBI/2kg6
c09YlIuByTBNPaOHUydogZ8jtb6QnRdJRaopehtKh6FNkjqz7RhESCCUxfy6wXl9
MBZ+1Hjmdc4YDoszOQPxV/AN+1ova8bk3R+bXwYnCtj1cYq0Y3G8lu4NcIgqHnj0
xR/sKsLbHki/GiXF7VocZ5sbqD6VfOOEEmJ3xDQc5j30ippVt+bY/VboclY6vQuG
1SGuE1qvcXy5r/bpLA+i4CajF8ce3kvxurL3l0U6DxAIrn4739P34ienfJzyJI9c
WnuyGyl1ldm7KGtmUAJSfCDE6Yt/EU6flW/fDo+eBXnqo1ZEBFQ3InNzGbBrBHRZ
ZYzo0Z4zalo12sFViDFUjKN41xa0Bu3hRoLJ/TMhoQM+o/QoJkYc0X3y9vx7K0ju
WCQzbr9wKuh3fek8Nk2h7tsuU9zNQnl8/zbF0WpKou8u7S6gRWtSKKdlc5MsXrOv
nQteZ+0e9fYPNqzCGFh6FaN8UaH+grGJSwwM8UElS/SU3tQZKPxjM8B7flcsdJ8W
vxNFC5l9pewFiIZiWKAPAQpZqYdPJbSbTZr6JmmTCeQElnvLZ+ghO4L4OJMe6JNG
+GdMED6PKQbErhY541MjR76YKN5NQCFq/Zf3QE+QUTGIW2/4+W45pBXTiP4BcfJw
dSXRjmF0ak4S+PF6QrVqqdrTgezOBnU2OvCQqbm+sGhFkzTUh1wRqLpx3bF6AO5N
RzcLlph6KOaRcu6LDP0LXZvXI9dmfH2hYnQSnygrpLo8W7FfL3xdYJA8dEhVh8XB
JsNKqHAI3x6EPPs6KvkkzaUydp9KUiMJJmbRlzT3tQhrM4dFs9Xuk9r2kyyi1/y6
azejJ9hqMF+OAVSq+1ETKuED92j3jkyHGo++1LkZc063P5b4Siqz1BUE5UIvU+bu
fIpI9m6RudswuTcNY7SEghfHlrz+II6HN8qNWNM8S8NWCOejSrMZMKc1hsm9NNN0
xiok031N65bBgVQ0zBeS/+01POIxiwJaVXUbsASyS5EjUoeo0nGC7eVkW2TprrFF
M8XvBQ3nyOPDr8pFyXZajn8WniwyclIas8kBR2dDHV5z3L8p8PSL0aKQweGcd4hf
BY8pHcObKbjTp8NVdnt7E7S+5ieeqC8hXO0Rw4fdYwjAwxuzHDoGiQfhGHE5cEa2
kzNf6kd4nKKPRWuLYxd7cvQ08xMdsvQksvdUrxn2MeNSyLsqVVyOKp76vDUSYalb
MlkWVF1HMiajn95MqFGR3sxowXxiV2E4sal51DJGkHn0GULzr0YIs91Ev/Pzv2Co
oFFj5TZFEc8Al5EfLPPZbXpclYBGBtPSTkZy2y/eWpHAzhfecz+6XSSAs2zAQ907
gZ+DkeF922X9ejP1ip0DGtgnB13Sb8rj4UvTLYfdZgDcnGf8jclGBHxGwRpaUyIQ
7SdmA7/Tw6VTsBc9kS1n4XtYwBH2OWB1H+w5d+QSCp/cHpMN1nlhSk3Kxm/oQgDI
uGhfg1iIIX0e20KBRVZ+YWy5OH3On4Og2OSPFETw+aVwivhTg0RWwcXBXGgF5H0W
A7qZ68khmpKAIDrh9FuCVVUrgz9ec/LXc3rUxYYylJ8VfQoVRJ0bL6bMbzpNEoED
H4nBaHcBje7aELAekKH9jJ0gv8VhBIaM9nJS0gfJxzGhXRyGGlX+5hoayPU6zLx7
TUY3deL496XZ+XdQc26xcma1VgnnqVx0Dqq88mfxp7t0umaZqgrcJWvwA+i5XRsW
3um+r8UuCzomp+s2kdYQKvY3vfic5yWuRR2e44q14yC8/Jr/ER+TOSk89yQetO1A
CoO5iLCoGytf29YqOPGa1kFiNjKjEb+Xdc0/lkTCgf90tEAkHrhcU1xeQ9qRuiFs
FJvXIkrWx1spo1RxHloOGcTpNxkmR2KNqJmVxuMH+t47xCuALO5vpWcAZN6gWimZ
W1gsBQuQOH6slo9lgPa119GX7N3wLhNCg1p7eOYuuHjSF0wDEOaM2QJl5un+ilAo
X78qCiUdbZ8uaqEczeQqirtBTfpPLly3kNg00G709B8HpUmcyHgHub18r3EQyozj
5GwXbXfQFnfEbXgQJE/njQq1rGmm2OIZa9Z9nswZx74UqqMtc8d6IImAPK+Z8gHL
FyA7raDUlXe75YVTiOT50CNLojkUclG/zS/YpOTYrlfdnL1Izqrs+pZr7PyhtcPc
BGL2b4KLUfJK3oOLiHIf55leNg++2pm9/CKS4P7mWp4cIESMyl739EXs0w3kqeB3
LuBD7jIK1E7PrCEVFBxtcfXuFXwAQ4PcUPp5FsVNlE0g/BMxfqPLnabz/NntCCnY
BkpO1tGFhFJLqapLFgaW+eGOiFC4BryPb5+f+AR81khPGgP+sNzWGIbSJ1APvOq3
DaPdoFPIdFoXmd6OSNuFrUm9/yPB2MNVeeMvRVcaEpoVKon4RclmWhaLnudJdV9p
igrY2it8rqNLvrcAEeLvRO0hkoiJBZgaFgK8nn4UUanZ1WECwsgZlZ5Yx8zTB+iw
UTOj4r+Ft1/nydzrAte5a+D4OuqeqcyBgzky+7oRnHJwYNbbhP2bXNAdqsOyIecz
IJPO1fXQDgxS8jxpOirwgphXbryPrgTh0d4XxEwbTJ7VgxQQPvJ/rPaDg9XB+Yq8
olCV8PlbtEutYfPbnNrKQPzjahz7RZjU5COCiUPGbrbGjra0E/p1kJDEC/YxpPNi
tybm5lw52qRJWSyeIU6x1YB4LMLcAhC9z4ewInPkJ9e4RBDJ+O8Iirpl3Xx+7awc
83pT1SngNv/fzHmDBvFKWo5KBnq6hNBrCirN90B03woCcB2pX+QCddyOAYVC+rnQ
xJzDflZp/aPNBVvSn4rCoEA7TmU6l9SJA1jXpv3Z90rPoKY5QXsAlDYmcaqQmSGW
/7o9YgCxNs4589+rk2hAD+8+2fFUDq4ZjGykeG5K3q/Z9KM0oLV+PPZc9yAf4umv
95uWncI4OzmNbeD7AL0yRD1tTY5wdj+3nt7AIVFHqXvEeVEfda+cKPrdZhO2/43n
hh0o7J5LmnXnvknyk03YNbrLDWpyZ1Yyv63cITKgzqqb8PMgX9jMFNwwQyQpU+Ts
fQ10jnU7rqOvD524NjZmg5fIY0ymW7dQ3WvCFZh5O+o2rJu9zIMvttjV1EFbC5CI
/mAlZUAvbLzPwZGE9B0jJm+wX3doSD5v8VGUc0GU/uTmT2LHD76OKasR1fAL+WEY
X4MZ6a5bXhbH5vM/k1tFRwVhfzr/Mvi51lZEEJzcoGosGRp4zU5Td/SLL+L7vW4z
XJQCvjkaD+hoS5ZxwYJbOngZW7IZghjMTHvU+bBnKbZl0h05UmSckjgCavkqcf+e
s59oqNrC8TyJ3BVZ9C5WRg+VIG6TA2uyhXh1/LQFYWSxASxv83PXeFGBS3Vz7SIu
+VwQ3n5W1QU3T5+Ao+AJ9FIdhq/DnHkNLPdAHl3sRMKe0khA8nWAH/vT86Vmb9L5
x/ktEAdJ/hX72h1sPq8KqNZHW5vMDPJv0vOCGW0miV2P9EnQa5J+pY3CDptOjsH1
HOpL5GArO8cCzvdoAy3sDi8+H/8FXCS4cVs/GQeVUQQfEQeRokkrLaPnhluym+Xy
HixvR9fk8Z3w4zdybN1pnRmGCxXijcs4DYJiJNks78eHikpR/cCGDFtyjlIdHPcW
PnK3mhmPcL31fXWnvk0JSVP7KthMv7I0uBNr6pGejj3MDjwUVr4jUpFxv3Hz6bgz
0CX4QzhKDo0V/6lG/U/Mr3C7AFqeY5ARQpoL2gKzlP4wTuaju8HeLVys81KT5u/f
e2HwgLGTqr+brAw7JFdRB0Nr1Z5+wCPLRsRYfbuF3GzlbxwVV/RLNxhanJDz36RZ
sRYGvqvhJ9hqOX1PhR7DuxTsns2GAwE1VHIIR/EmzAnM0+ZSBCTUIgZH4fup/ynL
V4QRj/2N24Wi7nZydA3nENfxb9hdTCTBhzYhZz9Z7tXyec1tBByIps9/5AxAU00z
O8Ua+QFhhwer6gjgUzDIEIgey6LOYzxA7yGh0tzShR4iLBIid1apddnRBWFFyDyf
ihRBH1S4HGSsXUGCt8Ne569Z0qQLhHHSKWJ5WhgFiuxsGcEFiVk8Pg+M2fEl1djC
Jjh4xrz1bhu0omNBIX+LUNPqLMzvwnNpZ+KpZ30DbLzKlhpFY32pn1H1mIjILTUN
ZkN+Iq5B0yfrFZB6LWYZbKHyAFQkw4Gfiml4Frrr2FPNqRleNknPfWW5w73AgiQc
nCeFZlQjNvRjbvun0kngF9bBIMOp9j4j2m+HMH0z5caTgLm7MobpWzMSLI48DWfJ
o4zq90Sgx87VFbRYOBIjIbHn/A0E50uNjleqMk733L+aGiyJ0S0gEHs6GSisH4oD
1o1rS18fmgQ+owJY8Xc1Cd0T9H2Q8xITPXCw5wTRa7vTWsntbO1/tNs4cyCMcEjn
x4oxDq8hoWdU1fWSHfG7Y4K0g3n0LR/T8zsr1n39U5tCcXu1xySF1ft4W/EqMZu6
IymzQWk555fDIarq4QlMfVGSFUNoXmHzawLWl+Ti0Q0+kY0I44tabHUvdDVlwPy5
r99eaN/4haIMCp5MXzDgfQ3PytHnEVlrYhCGTQfUNMuvyzh62Xlbf8hOgAwTQmId
Pvbhzq4brUL3GrLvY/9f4ILPF9S1s9zfYMHx9jSKh7/2xyD2UtN59jCUMkiWqzTz
wQvUAfFAbCR7muC5eFO/hwlNWSnh7rk3B/h/+L0CEkt7thV0AYJUoQSi5DZBZBZR
XQksi+fT5AfBX2X9r+FWm5I7f+dfH7Qte4xczYIYOoE3fMhyixP3YyjW3nv75M47
u6w1MlcmOB1IVVnw+9+nomzZr0ItmGdd4DmytcpEVGPECPfpfQpyV1L4q1E++Vo3
+eykIJnXWnF7Ywsipmhb4TOs1JMXqeRQvJlB2cMtslg+D9hhsh1BnXBOTvmDJh92
4vah/kNOhx/BLloUjO/4YLanTEgbGUD8vz/LXUGTTLNNFV0P9tJ5BKDaHGF5a8tx
knXUahGLCphuYVkGK3Ez1f6aohR6YTgme3ZJSx1+FqGrWZFwKlM+yNfsEwPIl1U2
t+lkMWisd4wN2IccmhyIU2u4YIoJFNWkvvhfLbcUxuOCq+2UbhLjLAZTvS4TS9v8
71mnlxvW6Xik8Mb9EF/AsDMTsu9Epll66czzc2fE/bMl02ZEin6fScfNAsMCSSVW
H/8N7KFy2YpYsQZxeAyXYx03zvQesoitvoldixBPUNE38hUd5vQu9CCBv/+R5kfH
1gettcad5RzHK/rTFQ9ZFewM5HvYIgORlmveaHSVj8o5/XnD6IIYV3dHbTq8gkjm
DoYLxCos1jGJLod234H6hrOlrfdy+vnp3t2xaZ0QJ7N9XSzKExvaOmHVQY8V58BL
4CS9Jk2Pl7pBEWcveaXZtc6GGWmWY6QMepLsoLsrF2bgi+9zBK6Th9tzkeoo/3ex
mJEAM//pd4wpmZize9vX5kVUPvxUehrNjfFc12VGop1P+w95SFLzOfolrKCxhGeC
RUKHFtn+D38fVijTF8tS280f7dHKVTgLW5uKLWAGueX8sCxs5wmLYCoFRupZKPrR
9+pwWubQOEL2YI/TLrkzZYaqHpxJqQPhUgy+AQg6kfcEiyBs9zNrXqzE6BPQtY+e
2fTr7S9GghviTO62mPU+dY4S37PVSuhhyLvrETKSHSbyvXCPGzwxUP08YMDvh9le
2yGF+0JsmFY8fOCRamCE7JQUcRnPompTV2IPvzjJd3+8cbyjkF2QyCxbEXdw4wP0
iyv/jotXqEOHCsxcgq18HoFQb19S1jxLa+sSkplDLt4dAcwL8h7igfQ5QWsQcgeO
l04EHclJ15qGcLsS7bxnd9bd/4TffAW6kxw12ptg5d377LPb4gblAjrajNIkP9k7
NVOlOZJL0dWr5OJw/HC9wzXPPbCmyVlxi1DtHsV5RZUu4G5IgVwADwdpZbCLSgET
OeznKImsaDq8iSaoCoQilvt1+J9fh6ZwyzW2c2eyOaukGdM6pTgzgZ3HeKFIt2w8
Ub1sb0LX3eitlteWHvZfaiZ8th5awsuxUawQ6El8VPUz/h1bbwOOCMxn9LGUUBF7
YxdMkXNIhjf+dXKlRlnTgYUmGuMQbcCXlKhM6DAdgmBy8rwV+ixJj/NG+pD6hHpI
Ufjdz2VUIXA/ojewi2YCpHu4lJCL4+C9zXM1QLE7Gc3woMR7M2wJW84SC6U/fAHK
hbYUUz8j8B+bfwoDNUqSiSWrvz7THL2pcqxCFxNt/Lx/C0+xgUtgHenBbB69U2+4
9WOyvFDuYGV9lp1vD/AFI5uFKkcgRpqNy2LcQ0HLDrV6l4q/MjLAqlLJ4Bn+AfuY
tdJcQEW6+ZQQ7q6oo6SmfsgenQfARP9i3Ww9vxxp2PiNm+Hhy0ZpZFD82XUyjdcG
S4D7KonnYlogkuE4/+H96qq54cm2OKeANe9+HiKvbqM0DaIHz/Kz9kx85QzJgyEM
drSUYTac1sHqpwjG416iLyz902B3KiXyrAsnuW8lBP5fueobhaf/wizh/ePll/by
1OzcTUfRtCLSraWTeMabyNIG6jj0NP1XaC5+nM9tvzWXN4POAiWNZeqrb719Tqa7
eq0K1WZKiuXqEX8S2+SWMRRA4t4XnLiHPHlu6iMUZHagWWaDUPVaqu4yAWWYCAkF
JQNUhbVNyzg8gH9zZCebYJKL2mZ1hr/GadHxDKGOgQLTh3O7+ogUS8l+0J4PBH+7
LV0HZj2aTRPgEKSLSZKtu025ws4utdTpKyUjI/+2BlwMeeX7m094i5tnVspVzown
Spn4nFHfxJJYo/McPwULbFXBY28EFfK4JhgOoGznCusZ257isRNutp3sQGAEiYKF
mx9bkiM/EcA9VYV6ELrUrBtOxtJknA5x2seaa9bhGwijVqchefyECJtGNMkurNE/
EG4OsKlb6IG4g9kXi1SujDCZ8Bm8cJZ101/FLGQ8LopWp4X6J5EnRVkoZfHkP65U
Sw3tDKxCG7e2nTNZ1FbhOWna6nwqGd4A6UvobtGDeJ3PHBtmVGNPIcWcdQtZPeP0
2wTNKhyk6XcmjLNiSQW5pcKwmRheTuZQLcdQLKVmY9rWgnXl5pH6X+5+7SD/SvDV
S0wZlKNRNNFfQcwaUI3X0WwJoAm7RuMq/MukWkfGVO5tCngz3A6vGXz3+CQXqXth
3kY8WuJbVFYzAB1S1ba3Tl3YSY7cDhNr9Auy7mW0UMNH+LlDY9ixosyvLCg0E4Fj
Ls/Bqx2y9gIGCgqXEZVYpLfAhBD6ZNt2GmFal6m+KBCb46i5bSJ/gPHQYXgl7yjd
em5TkimVuEFPrxkrbgvnzub4hVAH6r0da4F5v8fU5+qYN/Ot8X0po9CUrno3l+OG
11QWz9BMo7jwwA41nAWEXlR3Jrzc+8nnQinKLuPZbA9nB2M05HfPZLs36x6liudZ
G/+LRELuFXi7HebK0wVSSpfM4Jit8HbOncvayqfp1opyu/DMXzvm16/1fP8btjDs
fZB3YhJ6YzMLJATPDeamc3KoYmb3ZYhnyDCKC1wFTRxYPVd9ynTmzINgyQvzBVLB
+Uh5xr+0qqv9fh2xdPYSrIxvxVXoWQA8v8ggH7wMyg1i02TQ+lpCZ8e4Fg4rrSLB
kpqfmskg8AF+dKLB55IxIUjLPS3DTud7X5qS9CcFtr5tqvsdg+XDtsZ46cbuMzc3
oWYxEY704kSobsMeePC3bwjvhQGgSYUXlMxsOqPFzQdF8uSlA18E7pEnCBrFt0hP
H1uBwetNLjf4tce2KGu0RaaXpA4m7+IHOD26E7vTh8h5Fmc3ELd33zB6yLt4NHd4
fI7jrrpEKluIQTQEt67fEefGmd9bvHdw2PFtPiqyUn1XoSjLR1Sq+e/J0ASOZHPM
3l7gzrlhXeDjCwW7ZJLLrk4Low3fxETMds/ErD0n6iD/FXGA9FbuP/WYFj+G4a4V
47mxT+Jq84yf9VfSArzKlBBosi3WBpGkUsLrNpETZLZlDQeYlpXMzqHKFOUOMSs0
Y04TdLc2q1xJNGWJv7avmPLCdj/zBy6iliX5BdFxWnnSJ39rBh5gHnaAu1t9ouwN
kiiYgqfX2tTTucvynO58qt4zHCUOUTh7sxUQIWZ/mUHd1g5aSel65xnLs93ezt9Y
NJceqZZJDcbK9/lAB+hqtuV0x8DW0LpCfN7j2z8jIQubmCmvJLAGHlHgP8o46Dn7
Qb1FNLDyclgyq0Uhic+7w1Rj4FzDNN1PelsB+1sCO99jyeLexNEjzdgmV8JIsQL+
h0Pk+3lbWhG1rrbxAXEsp9LA6Pj2TD6kxG1wEU8H85QVwlkWvUy2fu7Vq1lz7z6U
QTEb6kFRbs4js/RMpVgQdKdr/tAxdyCjMphUlOPE+jq4wtldiHWin0LfAyEYG35K
YL5kSAd2ynNO8va01cnH8fES3SWsem4GZkAjFO40rVqBbp64yRTzvhOWnqCo9kQU
r31U6ymQWW8tUB0JqjvasKeTZKBjf0CDqohl7tYfF1lJ2XH+71aDh4hFC4XvLmVg
dNHjj1nBrUhJET1H5jkBoAokofRc/vbJ9Ar9OeB3JvRnGR9xjdZhLXbPenHDC4og
6QMNV0pOuxw2rGqw2Hc4zOF2hPVURr3djBx47TFD18Bf2LjKFM+kFwmpa9cUQlq5
FAPE04dFIG8fobSzVkZ//s1qFvT0z4hNRUsVWtiiBJr9+u/fIBmJMetrVxgw/O/e
a5tI7mFNTZASzKHKVcYcod/IvA3bb/b1dXZgNx4Hv2B+OSwxNFZ4rqyg0Wxi9UFt
MiyXBQD3YNHPtoXDQWMV2SMe/RhO79un4IsJhyyan3av4LEVTPA/E0fC+MDPQ+Bu
0Rl4zvxQVZn5NbdIOWoWzhmjE3LQ373Fqkmm2k1Op4oPyvYXZlA4cBeSKrU307FN
Np62K07akoohwBA+XtZs0OkxklpcX1CqglJYWPORg1lXGqHWWGO3VyPW8H3XVIHU
xAtu9zpelRKn3wggR3p7z878zTNwd7nHXSGSuo4WDzRDT7exJX55Hcos7mhBV0FR
39AXKynDWjoRQO/bAwY2RsrL4Dgkv/wvidOJzIcovF46DC1OBkX7mPme5Lhiq74d
m9kM0XsfEeTeNvr4OygcE7ViPkdlTLQwKQPhKT2GVXo2WPl7U60Rml01mYQmeq79
te6/hYOoKK2eLDx5OitYO9Ggo1mbqtaVZ7xIW0DX7UW4on/Z13RnKkI9qOY6uLVO
A+RY80XpjIKSd5xg9d3wQtAf/mNXYtGBl6IVVWxNhI9pHuGSoylnf77D/j6QIDua
yIT+FrBHMOM4M4u2cz6ws1hMNBug/JggzK6SslpfuF6Ba5UkdBW3YS/S3b3ltslb
sY4Ed/u1s0UHXyzLpDZ5HB3cznqRaK+nChFHB4VzJbypJ6tiMJhqdNjB3aB3hK6b
zKVsFXAkGaeiQjSm/xcqLhlz3Absq7ae7AsgZdmTZqUqIlh3t2hY0gxQhQn3unOQ
5t6RBNVcGfwKqPivg/sYIkGkhZJQraKO+2qctmlyQBH2xZRDMkiySl86wafhAHQq
1XHFLy9bMmmzPAl/8hQRb/mlmX3ZYISVuF7EgonjIss8hea3/t8zDGnrOviSmajR
vctdT1rURxTy7/qhr8phS7UTnAR8HTVrKXfVjHJOLdNPpf1SoEnRwVomqGLJwirb
WEd1sleu4LYsADGPdqHazT9x11WqcTwGyigUcHh+QKOQpV4S+enLuufAhFUfbG1Q
r2zM9ApvKtPE3oFwd/GHyhyQUMOK3taxo4ld1TwqMYxlzsskADOdMDdClpXlqR5t
cxQ1cZE++M7BkRFAsIjADHFbQXsP/sx4VlM0yaBhNKeefax+whxKvouv0S1RW/yr
V3iCm8lB7+CoP5uyEwZTDixIAjYAioEVZqncRafu/35rpdqo7hOxWSUGToTrXKjh
gycPUP0hOcr06f8bbkVyt2YTSJvtlNcBDqC4J+AODg1FQ83yyKf8zIuFUhIej0Yv
lEkOo06F6JlaOtszIrafZmT+iJwdpq4QaDRGEfELMFzfPdbRuzQz7FLRNxza2sMA
SWXEFpXlVrVKzLMkIndPGxQxRUIOxSqVpJwZPyJumfo4DtcTBkxu6+TcGeLGQwDn
vsx4SUSkrPy95Jcmggjp3a/oHVd9D6L+jVK1IFLfztj0tPrxwTRT7s6yFSH+EIO5
nzsWtuBiMW1F3cqu313UosNJvKbiFPMQLeKT4gFdlGiFBEZ/1EAX2xFarbxUnOML
kQPfj3xE/v0UtUV8pdspblrXwl3IX4C70KOxoxtJOJ0WdNTfXIz7OHGSX5sFXPl0
xQQ9CvGVkNeiSSNR2wJCVPZQ02cyRS50hiW/WHzPi+5rV2dBfwRfclkkvfJjPd2L
RTnbU1xdk9wp3fjGIRYXhbXSilxDFUmNXPZ/I++rk8PUDh+E5uYN04+7vE7QBL9T
Cwf2qxm3eJT68G+KjTPmUicYs7gQgW8A/W8gqF34wz/pb7yb/mgfycomcw3OfoNI
UABUqljNoFt5fHi0fkcZnsJm83+g20EyjqJA339oir4FO2fxl8ENIyqAqtOcnQOY
RcQxzpuvdCgPAAGav0/KeXcaiSqTfWNI4iV3CfS7YFEIxL6Ruct1i7AnZTZEIAbk
O7fJzIp+tHCYJAfUoiqy+ewOsbeKVXfRCo6bLZU01PjPzsCxR9yfrM+7SFMGVCcB
vsFDfRCNNhBT2zu4OSbjQ+iDL/u4cyafgvBp7fxETnrP6gWxEQJZ4VSG6iziowHk
uv6CBCOKUS6rM+9atLXAVM6ssPsz6O1cjzrNr+UffZEhN49o+Ci4T2W+Nzm2ho7b
ZkuWr+u7epgIXbwfQCKPe/6jiFzgnGgd9Cx7KLJ7IoXAMkPgGmYpOXEPq1soxPYK
vB2JWI0AhnNHvmtCn3C4SOkbU8jBZVisgfCyyFGyy4GE1jTZ4nivJXG6jEVwM2F6
4Ecv+m3YhABV4ddOt38ZCKV/GLZjxA2pDMQ+FiIebrznH4GAX+VmMPd3t8fRHeXU
UaOYhbcUCQ8LP9UD9nXLoHGLs2n6APK0cVABZjtOKxdALWzWeRzh7ikvsA35UHwt
b5f5HeHCd+PSC6pRbDlZ5Tl5vHjLzMGNot47g18AbGUalpq/LPjwl2ZsOFpOPxh8
H6wvwmzwAoSj6QvwXHV3dugWQt8KyrYIQ9OPpNdo4tD+Dv6iMDwO5hUp5SYMNAuX
YxGnU1iTlkYlZVZiGDT82v7gGUidJSpG0ewp279+X82VgmFH1LaYEwS27KfRIito
VI493NvpL1MBEo31fCAUxyAUDSRoWGVi/9UOLv6mlbi+IJ67Wotme6whvQbCAGJo
m704Fg916gdbfgd0uJOLggA/2twRFlAnqDeUHMco69gByupmRsF39gy9/LNebCKM
4jw5LueyKwiY2KH3TY2ILoeQDqnd9kVfFgOpPvo+p/z9/6lipJ98UB3u80ynb0Fs
3Cd/61rOVjQQVV2vjbZmGnEAa0GoxRukdMiqZS6Cr4xPAfZpfc8hfVuyuqtjIKsY
BQ7BnUuukUulJX0pUXpwS9LSEWGGYtQGOe8EUlhRnq3z4lB+6v7zXOdy58eqT0QJ
nfrUBadivZpWZiI7kgEoc6KjkhDDt56GEF4vwvPJLug6/lj9kRY9RRaZqNYAge0T
+3wDWAdYrOlLK/GcNXd8Njs9Qe7WZifEfXya87epyYI6cFSpu6ZwK1wJlltyDR/X
YPx3q0Z0175TOPo8RCR6h3L5SFMmxi0aKE0jvIeDv/MRHZO0cswajgNP8+XV3GCe
uBESgGLWZ9x2NkLhz7XWWJK2dpGpQI+rsGdztRaTXPshUp0f5xCa8UfED0PHAWzP
sqljIIzgOtLh5vDzy2PW5w2BpjFVeg7KD+jgKh8Ztf6tDsiQEeCikeT5DnfpgeeG
dwWmOU9/Nma3Zn9Og+6+K5Ke4LcLa1gEmHvFnOhP2sVnjY+/lb8nUM2132/cKpUY
XaT8R/lpHGQEEHOHwUcFPouVU4ht/uP8YlG7nOxPgnrRVM7bjT1ohXIzBR5UCVCg
0GwQivrxgWpz9XEfEZxe7zsiVCnUExmTIYpjj2b/9qvjUWq4KsQ62bQwos+IrcLm
N7Ecjajw1kZub8g0qbRg9L9erGa686RrNJwOA4TkbWh628EIab8A9JoJhzfKOjTR
ZoFtS9UXIHasNB02vvd/NKQEy0G6qAQBMhqf0+F/9yVXvWL+w8kW0OudwHrs3xUF
3h68miDwZEmuuWEi5YEv/TuChqW7fNO9HN9ok/Ip9Tl3RY0S0swZdbwvJum+E0GY
Nl080kuyRLKhekexefs2EJ7n6kk9O1PwajAl91uoKw5WKI2UDO8TCHMnXYTRD3wh
O1jK6EG3ljskjWrfHQGVcaxPS8B3HvUZ0v5mB6jbjrx8LjGgbTzwUVIq6hG9i8v5
i4bBqYJ/YzRXW++BjTyQX6k9OhB0EjToCZA565gSA4RqFkGYNFDSx8opZ21xT2CW
x7zbsPd5Op9qM2KF/4sjlvLgnLhg48689CfLNLpd5qGwwjt4rb/KCNo+ojsZtFb8
67Gv4i3RsXCw5/Js+vnOctZZ44HiDLVvPnS6RRS8LbOLYVdoZctRenGhPV80O4Cg
8lo6h76f2k3QUqC+/Am/LPKRiByplPc7+eoY00RsWMltHx3EnuZeZfTngLxwazYL
utQh3PwMZgrtRN9lDfqWbZzrVlYcSB6zTeLND/fCZoMynNi9h+Yvjq6uz6De/KJK
04iv/w92hw9vGc5pG2fToOklhDfVkQaUi9ngGx9txsJ59TtEDsRDC+suNB/37V1y
5ddky6OqeOPhpG/3I8PyavSZlo5vTgjQi6HuLriNvmKcDcMdo+Ug1OVXidk2TJW3
FWi6ZhhHaeYHQ6+ApC/D4hxb6dIIzNqVj1ji9r+oBH/bvLSHpzuULA9jWCyigRKy
wY01ZOFEA+KaUvh8QUM/AycSm7x5qR2FdbWmG2G17qEwTBHSJoPUCrdUlTIh9Qhv
jSI4245Kf68ZQHov2HUbtlbOpTvubvGvmEBteVD0/nicbhIWComFkb0lqfYcnSyS
UM7poMVMA8tJzzvfBt2Tst5najTV9DcwV3UUFVqeyFipPEO+zi8IvrR3eQuzavyo
C1OwHBbSirJotpidndT0djd20am8mFu2nSeEDeNxO7m9Cva2cQMGsOirvF9GU8jf
8Wmw2mkioiSVpu94WS1aDxqlNPOCnTXzt5rXlwDHNh7YUT3LTmiQSmrR+UEKuNvJ
TfG/D3TA2HTHvPch5Gtw9wHmQ2Q2JcfcTmtGhNA4a3R2KxAjL6ooehppHBNrmksu
kZ6aeuar7JpDsMwbFBsfZ9X7NW8YfB8HuJSiaoMiVV/PoOWtjahZGzYWR14L827h
IKNvjdVSbkuD7/LLYzCW84cwbj4hnAoL0Rb6Nsb5dUVVlf1E7mKlzIx68ZG7DtXs
3govw8c45VCRW/AdLl0x6hyipRnFrXuhhfJI6MZkoG7Qym0sGIO0gu0PdN3vShee
rXXcjpxHB1HDthxgjS3boFftYZe22k8bE02jcqbji0cx55N9h2mHZG6mge06aX2+
LQLZV4JDOJHeFNWnzAP1GAAE08ggky1LuR6DEeMdbFbfuP63ieDKtP+BvfJzuuyS
GKl/nCjGTYOuZVdge6ExrNLRtmb8ndI7tl3UbgCTYadq0wB2IKR5fAOXf/9p/Gr6
omU7xWT2J1TFsjfzAt9rAmHrfILix7xnija4UCziILyztoqkWQrRPYmikixoKRk7
tEDxZVIt8RkvEuOoMNTUGxMMQwELCXzSo7cUEnWH2+1+M3r3LiTlvJK12q/A8L3d
O11izwxS0WulR/uHwuXYoc2kflH3P4vpcoo9gSPbqwmC/TEfg6DqPd2CQAHB2fO8
WLj9ZVBfqCsXpGh/LGPiezbNl8O+D6lQYamSpXuVWk3ZNS+r8dBXIIByb3sMTl7W
5PBl1jPCwxD/AI1fYFhp+SReG6MIhVHDCAlaSmrN9vec6S/i7wKzkMF4LsSvhW4z
R2PlIBRf3kM8ZYDbIA5lRl29xjR07pKRYQkEvxOOyxtLzIGNIfrBYwG8WOl0OXXI
VsXcODYiikHrAP14TK3iBPbLp9EFCJX6GEfS1g9J/+xuOt9b0lHzUVDTubh/l1zd
BY6GrBDHLvhVer7V6JWwyuGU2urAVDpNB+a730kr9f3mXWgpwvONb/rsnNCr0AQ2
3Q/WdYg4F3XBEzIKMqOAM31UAFbBq5j7ax+4I2hlNyMnIZZY6OKYlSo1izpkWwbr
OSOmHEywOCK9/d9HsOT4n2u8rcguKxoRQMuZNOZzNlg18rqg+ioSI4oDgtllarEX
HKgjGAZGc/5ldGYCfGJHaxtXssebr0umc/U0e0CjxMsMusiESS61dbUwvtTMbqqh
AOU0OdgGmjE8GqVDRKM0iKnIk6n/V8v49h+rZ4kyWDInkPcX/45bfO3TSStejWui
/pYPaNws520LbGJndxUgR0KrbuTrDuDpEnkZsozR3Yx2iWnbygv8ylLFXS2QYVBi
Iv2PcxzBzIwsj3M+wKG1LHitcroA4LYz/L4j8G4NYtxOuqLx+Qh8/b888SBGeFLi
4xW8YqmpqCgKrSja6zMkkq5Oq7xFqbN85M/jWhK/dh1rmEVuFDxjT6Tq5+gl8qfv
pcae8asXLgPtFBTJ3cPAGjb7lcHANmq3m0mM1iQLN6ncyePgQg4XPexQTh4IUzQl
iH3Wor1USdp2+3KkVQ4HYX5ScLbc7/omS2XytKyICVO53vqeHj5tkzamjbMuxzsD
VA8u3IOQ+EbRYtFD4xOsjjRQsz5u+YwnAPS+sfjb4dHW0tv3G57zKo+TE9fUnrUl
iRIWqZ1Ol/T+8u/gRdG1tq8IkNM5kFudWiFZ/uBCvahonwU7zzELb4c/LcnsjDDz
iA+Wx85Nb9cCqfjNMIW4X+d2o/DWU33mediJ3DEdgdgeicxzsoTRssIMYgTikkxx
Hzwp8LtrbvbxXUrNznSddSRfOfEvjpz2qEkO+cVQwWtSJwSF4OurvHy47MIIeD5X
OmxJEBbxcc2WmV1M62VsC4zEaGNIzV/dO8uoxhWqArYd+9Tv0KBCKB4oRBbbscuQ
oNKKzcnYNx5s5Q5k3aFfK1wld3zjYZNtynkfrfBsRxkyv26OVEIh33l79BAYcI0f
5ZZnx0ZnuBs5q63KgHmFvbMRv/BX6mRIR5o3dHjlm1EdnrQohzx1/wQAstbP0l7C
ZQbjVXZFfWYYx+zqFynu/TUran83dyGJFiN7HD7nUqGP/Q9MqlJJyNhYl9aM812u
/Z+WJtmPe/ENddFoG24fxxYr48GGDaEbv/wB4PSGgGIYYSYVxDi9RGmRFO5p95OQ
MAPM0qSKZ6Y14+KSVTmFuIosEnGRzO5btqZQlOZAdwdPFZvwJz4FArsESl09jSJX
j2lA4ovFaT/Sfl1WbXtXkEeAgYespcr5HLO3nAfdv8l16wZjTruOmvKquA3NZk0F
Eu9rhkPcLiBwr6iBaN5Sol6O5bbegPtPobvVamTGXnuZjnUgo4DM0bSOvwjtWfrt
8swuAWmmY36amwKQsCykaP7g9mPcl21yu1q7K15NRpGPlFekydTMoPqJTDT3v30C
gmSoVVmWqGjex3UoZ1nomYjh9E/cNEmCn+drT8xzw5d0MCL/d+O6JpkZJwLN4cEb
0d1EFug4v2EYgL0rHXazDcYAnLQMRfhd5SfSKH663lcYXe42xSU/qwaN4h7AyeT6
MtPdX5fsIUUC9kIClhWZXIFhmB8dma/COW88R+RxaEoKOn+PLjuY0JDfBvjfMpaQ
LtCvib2LwkT1aQy8s5MlRI2UoURdjJN4o/nmCWv2HX8Xhv2w1mZL7uxYZamtDjK0
8CQrgxzve4dyar002K6sbPIW2NIwxoE9UwQani/lw1nv3fb/9p1buEkytv1T9oLu
ExPKRXWpSAR/eKb7Yop4fA2WlgpU7IJlb+sWQXPYviWMV8H8rZArpeEq/jWg3hhH
bhXyxScAvISJg2e6IR5hbMrqvOBI/Y8PdCrU1S0pkPZEF7tRVp9cnH67txJlD1iL
r9CmT5/aW+f/K8mfEn3LVVJjbgEevtHDfKCuOIbsZGl2O6e1TtZn5dxlKGM9/mdO
yZmgJMt7LsBa7WBtnpBEr3ets1t5klUxbgF8q3DI0ua687V40vKyeHbgGwln9czr
anUvd1bUFuQMdTL1R2+vMI2iFa/8TUv12ZhcMWV6qTRV5LPj/Xq5Behn4KbM4roj
75uybofM2BIz56D4UA8YdrlBzNbSWiCkAxtRrZ6jYk9eoGSiyDDKNSdICb4qrky3
q5YUrMBgs63EiCux2pKovOMflpUr34dPiaIVJXkGi9jQvsq2LBO+71Q/0YOozYm2
v+G/+EedZaz0xOVHVusyI4v4CWhr8aBmIBOR7wWcsZg8hHlq1qOoz9O8eyFMKWey
YcCP2Pmo7qNppQXlfo0N3HNFNZJSalJaz5qeE1NGM3AN3Uzz5clKvQcNdFAp2wdf
sIRSGdxp0v9vFneN66cgEqT56CYfTSxNOocVqi833M6PBv1Qk4M0ZiXo8nmxduH6
XybSJtyrxsOIlnWvLQt6/2CGyt7YTIiUGWJ6VxDb6HTh+K0P4zoJlD7EL6QFfyQ1
x1s4N3VsqsZTT1iGoI6mNBMRtW6sTIb6OivvwLcSeZRtt1UaDbh8A5oKgEA6szIK
NFinwOcC8ojpXtgqtqOFkTvcvGD1SlVZ5CMYHjN3nLqRML9bO9sJKe7zjan5mFyv
8f+O5Y3GyzS4hfcoqmwZQVzAfhWMqc2VPavHQAGGlkxzFt6aQ4S237WEO/CoQdpd
zozCHgfWsKj/rmlOSMgHGO8JHLE/6XtOOvkW0Ur7ZD5KXQYp4LW1/4BYh1EOcy/q
fSQ8ZY1p2ZyKy7xu0Rq3HLErw60SkEGvpmOwEug94VPAnJ8GohMVuj2Y5gUsRopK
wxGOPf/UduszERutKW7dCZVNge8weGnk7seDQpiufUWOxiKep4XZ1NddL9SbvrbQ
/smL4IwHVeAHJs+rtoYTZ4mrHQHi+CgJZe3Y0XQNTXnOgAOJy0Cxx4JCb7Oq7ole
AB2n8Z33nP8Toy+F3bru37zU18bHQXe1zNnYDbTKbdMOHBXFvmYxZVuH5M1piY7h
oZoun2y8JT49RULmoB+Yt1ZXLb0W1EXK0yB9132kVmVOBS0UtW6OH5+Is1vUiazF
xHe4D2+qHWVLNVcbkOdVLO5GfYlLojhAoOeV/Fyc9PrprnkhaM0ZWmBiNF1KlMsx
VyRtZ8VAZ81147OwcTwUaRiedgufay1/2sDBz/UQ/XS4eWVERatZi5mJWUTG7Ykp
BEA0f64NjC2fIE52Xdrz0wK3Za3F0kjhNUYCuWPtUE69PtTt21RJdN1JiLwUjvuL
dAIo+ye0XzL2Qvmfy/REn+l6s97wXjVSmAtO8lCUKMu1qhr2QocTupSNEzhFpr1T
+InXrMQJ+POwKaqrejPRmAzHBr55O2QqIN3ryOPyHhWASXLwVTYhlECTFGhL6B5b
tdMi9dqz5rC3V05e5zWUvNyNrmATcbHxpamiRqscwR40E6QYczPDBG4nVlg/qebl
mipIpGHuKX34u4O5i9pAZLL1C0ATji5GiM8RE5rVIWWKBlQlOHXG/hf6h2+EJVCO
WIjh5aga+hphky53YQuwLtKn249/k08jQzcBnWCFoKHsxRZ2z/v86CVHKGSKS30q
nf/WjQbJYgNLIHab1CjoJ8tfc2fAR17w5kHcEZ2z9Mst43fvQWRC6rnMk/DdgZUq
sdchknEhjAcOj0vxaEBHGpoSvWYn7ZF0SgO6yv3QuPsMC1GOcyaZkYYGjt/baOQk
9Kb2V/vq3gUc+0uVLWiVkAipfGk7Att5IUkbigkpTd9wEXiSQn/Mljbzy1HMWwx7
KLc5TEoAh7qZ4TjXM6lYjwH4uRYg0DwOAFwB7INC7LVX0U3Grb8xl1Ph3A2UOlmA
wJNpC7g7ytfcWS4wdUHsCXOsBuQP9y4sN9KeWPFMen9KglYDL/Jn3fPrg1PfVj6/
sAavTNR8HRaZWcMrRaeZBGH7V+TjyzhxwdVwYkygsH0HwHd4iI3fQKBT+47IeSWy
OHitDsfRjtqqea8E7UswxEZLKjDFtbBNAgIFQxBuHZSXFM4VGxixp3gRyLfg/WTA
jXsXCxbHkW4p068TRO70f+E5cXyA8ggxB4fYeNll0CrMic0CXkRlqWb4o1Wm5Hco
hc6Sh/d8TmXZ3kNVZ5vAyKIS/wBxYKyBUs8/n49fYtG8SiT9G646dDZ17aO82iSx
YSbn7pT8GHf5XRCgIpNl5onCWl2wY48PWhTrAO5Z0BfA/sLtIvDGnrybJkyZCQg5
SrHfl/mhzHebNhdFx5TRv8NRw6BKHGSPVkJR1cbmRbJkpHGBMYlhgKGa91v4gGNF
6/nckl5aFSoQRdgTn40BQEsC2gDJRk5HcWlhfjkMfTUk1JR8iLVINeqGb7PYdAke
btJUdlJYcGXYUzCvKz5J5A5rxX9UJyyKgS7N8LK1+RU/wAlOy3Iia0edXnz45P/4
D2PZufYRuS2AjzI6JhMWXHvhb05Gyekr33QVleScCNtXCPpBoiLHyN1go1JmxUsE
vjnntYlrlT2TVK4W8T6cIks4SMn7+3x9nW3B0NHtE704LlCvpnP4h7f9reTkeWZz
Lll2+5D3mBNiPU39zUNHnQ+mm8ok92sdFNgaKeiuQm4T+8IPeT/CaHeby4xkck4e
4UxrWXrA4XB7fdv5d6tOBRvc1aBUfbTiS4+QGTeE9nWG/VxQdUREvJe1iZ0BUP6P
8Z38KwU+wtaZU32AUiIGs4tNjTm5tbhl3nm/1W402cnF1u9NNn9xI8wLUvWYKvwx
b2ffT+kiD6oc/CFPYaMfhX/OG0w3pd6y1sWKnY5I23VuWcGSXkm0kfZWCagbgxlY
DKEaoJcvA2NImhebQiJ7P7UDKvC8OJbdZW4fcsK5WbLcOoD8/tRdk6ru1l+Mu7GD
i+z/ePfREZhnxUkqIYsMbNtjEIJ8eg6+RtKeXCYXt1r150aq28RZ2Pd+byGgCGlw
b82K+L532TGAXomjq9URCX7hMixa1GcvUPWDSnQRuWkox4HTbkbgwjxciKOIKrHk
HkBzRkxiznL104XZKooz3DOF7ar7vGsXaBPPHn/Mz4t9BOQQnWph/igUiaLHuyR8
P9+YcAM4/WWZYu0jXvKKOMThtZhYCDJe1X1qDk2Ni2ItEHlxQqGnMjjcIM21sqfN
nbNvFhSb459BvYnsINxwnT5waVqDhopDlRfYXkI6WsK5vuFZs9pzQQoFcbE6vmy1
sP/n2UAaU+hfFtVCQ8n4L4imUaIvViVxkvDSSE0e/A+mPxlZXTnVrdtTKBdMRDeQ
1Y+f/CWfjJyZLqpq6MiWlXI1rXjMKwJmVPT1zqgraNGa+PGeEvBiKL2TLxVzHm8S
XFcfRdqjve1cdZNDmDUPc4LnioH1n5G79ptLF8bCDlqU50FX7xA9LFtYAbKj7r6N
OvfZ//GbW26c49sSdSxVZuqzQ5Ont0VRxdXooLi19gilcPsD/pyZoz8Z1Zan4axy
2uSPLLhE88SM1WeMmmp7dzTFfcJPtAj0gcuLUvWHv8bUbREb5fGnouxsw5ELH5NX
mA7kA7+qe14JTAVOZdFVNbzPPhxOyJAvGJ1Idhf1yY3Q5j58Q7I8EoC3lwePhs+i
B2d33MYZ+6Bg5TpZulwSMYhOaoXJcE+3IvuGHS4fhT5GIgnvUJD/XFqAjm0Pnqmk
dW7n4pSDyalBuvS8zRUYHPUN6xlmI2SOU1unf45f8hwVjtjJzAJFiYVQVWgk/b7q
7iFCC7bHhl5wMui80iTbu84NFSHFVQ8hoK2S2ZTbCAFrg3KL4ZOyopDnfPHAkQ1/
CINbGhsHs+2rVLub7zoGgXpBK0DnKRncdIkSVDos1TKtKkkVhAWLbR80dAX3yJrs
AWTi1nmtK3gFuzaRE1vZBKjA25I2DiCs0QGdG0iL0WKu9dNEzBeUmiopv4SS/qJf
5HDX57KDLAFAID646+Z24WB1jrHbv3eRJ0AlCKCagDgRvWanwo58Zw6LyfvdO6eJ
IIYb9ERclJFUxFrSOidoBgS6ltm1wNH1otX30VjnR6Z/xgpWxHM061A1p3emXknh
GFVJJOABZtBbg1CNU/4eC8F2GLu0lH/tlmuNUKf6OY/rhC2o6/eqNzMgK7VxyCCJ
z0czdD1D3GAx+qfQSFDP+xmkz7kfhQySU6kZ4/kQL8iS+McreBzi6Nfg1z/apGWE
8W0gSfgPwodHJalz6SyUqwObKZtFi1Cgb+PkBXacCwuPgjyQVqNJHsg1jfiLEg16
MbW3gBi4nWA+HC7+4q6VVd2xhW/Xgt4NxgX+RB7kigTqKeRyJgubJB9ZPuHW4Qy3
91sAPjXkOwurAQ7w1WxTaBvPYtHoQ3GeTMO1iZEkCTKhYZ+CySm6Dy1Ov/lPS+Ax
8wak0O3lOExp/20QEeuci14GBnHe4V2xwFRGewUNv+E2rwZn/1XU/28X7XqBmux3
3m3dfzPsi9gtUGq/IdHjPp8HflU2MUWmZhnKOyZOwngsRCVAXW43yV1H6S78kK1E
1szwg2g68xi6RzVtjLO4KzLUWvIpr1QstplVWUjzxwg/ne6b4IM9HqIG7C/bdV0k
A7ng89XDME8q2SmzEq1qw0gWcK2epu1Kl9OeR+eBpobzsFPwMnPwb3XQDw4ZYcN/
m5aS93mT1Kw6builRRogWvuZUgXU0xOtRjwNlw8Pl4crltRDqGgWiGOuZ7nYXWfk
OSx1+3jbLuUwIHXQgkxovi5aEMDL1n9cURxg+rhbiznqZdi5roXEGAWLxF7d+TR7
otL9ch0TtUX6HifwdlnNJ+d/Z+wAI6r/cDaTFt8W3AB3S+ilKSiDaNtiFYBTnpyz
PXl1L8E3+zACneui3LL/0Rb4VTuoV/yffbBTHgGWCn90nZ9Z30UX7qZ/CnWIwhV+
0bKWpbLTkmPUu+CETusre+XLm3MhHgKuz2BoCqcx5oBcsqNb1v1F4FLNkIXSdfSd
PX3JUB1QqA4JCSG4R/MFVCZr1o/fyRPjVNEGu2DmvpyDhkb3sFwypPaPSVo48AAu
DKXzkoWEiDo2UtLhvY+M25sKVGuiICZQngAW35ZmJJyhMmVYU76fSAfsLbYmh6x7
MNY0/5bznC9IUOm+8t5y29B6oK9loDPh6Nhw98wCEQmoFQNfiqMxKhZOJadMUNqe
WDw8ob/Viuzlvbi9zgtJcPMspTY/gWJMFuw4e4jUMIkhMyQLHVNlErFapDyFIUf+
1Flhzu65DrIjVJa1Bft3ZpB0zJfLCAPCfLRzdHpEXBQitwsz3Kg1Yd3kXJ0GnRPg
F/Psn0AaIV/XuavQii7mOKx6RkWZvciMpYkSSeg/ZVZR+XVeJnDQSJ4c9OCJzuvw
uOjwQwwdakYG1ZmO0LI7f3K6KEYzc+7czqS+V5SfQDD2Z8DwkZvHmD7wxQ4w1OkN
cQq/uEIXZilGSiUIw7TqeUe5pi8xPM8XhbEIq4sxmf2lMoU4YZ6KoR8SzA4Pt5nq
gbkha7yEtsZuYu+aOG0XSD8C4OHQLjguW6ynOl6B9MAIfE+lGuWBphyCWqRhQ1N2
B4ADQmuetJf73h2DaSy+rTkdiaW9jjrtlE5kQnNOZb9/thnQgZ04nW5I2Ykp6sEk
frYqg/8OFrMXqM45rH0TQ9F3HleFgp6Q3THOVXiGcg89sHU7FUnIo0BwL/s8bRR7
XwqziWtQJZHkqWlBCgreLy78+0PsQ0eYKZxQqwBYAbrB1ozabv/XVIfptuihbjzt
ytlDQLjpD9C9FcS54NlkXbj0A5Z6VYhoHJkS460s9jSPKrvmEJ29ZZMEhHx2DqQQ
whhMcnhNfCvY5ktYIamPAdxPYPUmASmdQ0O86ymaScWG5T9zMAV+jtez3Jk25eXY
TeuWJO8FDfXMZowqERr4M+rztXET+jwvJwelW2pZY+cR3WfvqLGfKSqTNLUUg7wo
HI49sQc9+CL6IDvs2A1P0Xc0ALfSjZ92ucAb5gUR+yhS7eeszsCoq+Bdn+kZueVR
qj3rvbNLtJ4IxTIxn5yraNdm71MXa87nAvwUYsy39WfUiaFqaKxvXq7y5uB3vHSs
uArywStiMMokjZLOxrmSgvyBPlWQnaR7IZiHtyzUsjA4B/DOk+WemQI7SBciyP2/
diKE6b7bicsQUW6IAwHzn9LuGNF0FArwQDNHT+QKYa0PXngGjb9XiMhGjmiYtIfT
nT3PRhCd8jX+JysvD0MwDvzaChRObaZp5ylXNXQQr2DBLNr1OJl/Ngxa84my9PCf
1S34S+cKJSCdYrGJhTFzN1SW/EFAygfeDaWWRn+akln34wbKnXu0EHAWsirbEBcU
5jGhALmMmKdzW+un/CfIgyCO3f7Y+UwyCo3c6nVOEUgS3syvbKHTGytNp05e5Al+
F+2nKWh/SRYxAgQHB9HCro8V5O5XdPj3+kaGUchClzYCB2agE+TsWGVFMo1INko9
VMszpnFUL2v2t+p4RefAq+nmcaigIG/YOMPPtm2bdoF2sqqebeWxwdEI24hH1u3F
mxGbq79T4vQmOpOJRyFI2MKTP6kmK53tgmNLCd9Y63kU0KYH27XzR7zoK7VMNPcK
02QfJOXWKcTbXqpxMhBDvsINJYCvHkcEdclacgF2j7bPBIkNlh1qKE57qsagPIwt
Bf8Ci6zuhDGGUTgQvMdxkHHouuQNaXo3TIl4dye9CS6O+dru9CQa3A6Rl4pZmYhZ
sf0UN52GSswOlsOEmcIi7PXd7XD3LSfesr8wgzFp6jE2ncR51cBRIAfIYDm8FBgY
P0n+y2hufhoY9Vo2/iBeV8HSEyIW81/kqIQJmXuTC6d3OsJKdWjm/B+yRQUwYPt1
id6ObJticaXJVNylJBZ4uT7vsqJKNqrC3qCK/sPKn8Jb2mdJIY5C8WndoLXZwQzd
Ic3/mePKmBYTa+vwAakFi6g/VRsDzb/x5ezONRSFjNqt7ySB3O9baAMnFTgqfayo
hmA8h6w6zGAgwSPALdotlx0xCuwx8X7pPQChJL6Dl00fMY7APp+Nb8YP5Pf5cFdL
/A2HLC09I6HHtOmWVFM/aTu3PyieNdj9pti8PrjuMDsxp9xNvUtm1EJQV4QoJ9CG
Siw8jgHT+Wv6apO7WTYHBYMIxQ8J+9/7AxQ8hW4jfbRdhnjdhHyzfg6vr5bbSYcX
p0clWi0/RJGjpMkcgyozeCdalnu0PFLYRUhyWm80eoO+dPZjB/TWgRjPI/Q26KLT
II2h2smghiw5V7AGAo2wr8pk029oz7icF8UI8HBs1+/FRsnwvwLGVG0C5YrlU86B
XBg0DIT/Wx7IemZOiNTpz/rL5cj/lCl+L9seZHUrbFwH+iUCFn/MrdFxpbwVroZ6
osy/Kye6pezC2M8i+z2UOYVZlNmJYNjS0OzFnBEZKjXHEvdu7iqBGxpwl8N3z5tR
bEkRKsNJY+cm94JEHblslsigmzIosOiQq/kSl3WED4Psrbp5ttTSz607GuxiFO95
yiZqIzqfotdiHERyGYrSvmOxP4BU6Je4VBid24+BKBnuDSpBfdcDsyiTIkVfKofF
0IZBr/GUSyGIVXkzARi5JPcs7y/ZHJ28XsQq/n2FT5K8xk4sElx7tk4DRxGZGFwz
huG52N3a5Uq6TuofNRgVHWTeHSb/dWFCe8Ea2Y0xTXGecWK8dweU86IUad0403wd
CYw+b6KaCeEYEv6N8NrhnVhWhoRxxMiBQCV5b80uytBVX6AffrRGfE/JDs1TOo6i
4uANAFpHbQ+KFisTFoxfrpeWOKEitO6eFKtX9pGna+XURWCK6/CbFSDyfaeaEo1V
XvgPA/ASTVIkVphl3hOPE0JZBRBIAynSTe/GQarHpPXyY82R66M64XGYr4U3bjqJ
swRx/0+w/aT8v66/5ty61SICp45wGfuFIuLXO+6U03YUJjcvAGM0zi3xAs5zQQ2Z
YeuVleEM3RjudYi6c1Ea+GUlpUJTd6p7pbx/w5gqGpENP9kZM7RkLE3ZccKfhT6/
aEyS/J1cz8HhHqIBHG1C2OJCV7eu7R657mrFgQg1QuUSeInmZE8ucJF95nOS8jqf
pF6lMLzED4iGjqirDTliC0qU7NjDmEIAs8i1cmIutM1qh3V0RhFSVs5jLb+Xgp11
tfMRJA0a8ZfXAb9ObDKhqwIczjruOqppLnEug3MWKrczxygFbf6A/NUgdwxIxcKF
lIqmjCfw/HzmMt5zLR1DmupO2A4iyfYHgN/JqeOr0ebvm+JFcX530wi1GFh6BoIK
PzC/uqSEA+LagpPc6lf7xLNE36BqQaiV9S1PLlWzoOowQNPXXGk744ttmHRs/ZSs
eYCb1Q2B5JaHgsIAfOYWBFg//LCZfMWfW6Nap2zk09MCa7eU4ukxo4+2KOBl5K7b
ff8oIw6JfOP4wjVimbtQAYsQhdNoobpgBww8Ii++4j5KPExhNDZcLi2rL9XIHiyp
E3OAW9CQQPvTIOM2ozatAmdi8L0WxmfIUGKc1RSCTOdDBo0ezd0MwbFnaQR4INRa
BR0PwygJo5NJ5FZPHYHYEtAlSIrYEuVPoSNp7dzX5d90SQtocWY7NtXAGvWfh/Y7
VBpH5yxZOEMlNk+k8ftuLeqgKE62qEa8M4dQ08luVi9gDD7ADgisYWlIViQuyhRw
E5BkvSSJ0+8cl8nu69NLry4JicdTMT3XkXojj7LR/c4gmeXqtJFmxCZc4njJ+2tM
eBGY4evRqNzCmkxuFNimqH8akJoC5mDUKp5dZ962ZTtOuiVbDyeoNFh8MSFsR+37
1jD3EynYimIWFNpZ1NQEPQux8M3bHywHvhTrXTts2D1nr9z3B5yHmsICiHd1Dmhw
L0Xg/PG2SCI0/vjcXUt5pjeaOeGTjv/tu9mGvfWo8UPhyIOBNlJLyAUTL3Pe+6zU
AEL7jik+8D6aTC7Sjit0IxVw3a5yRM4TIJitKQluUpRNB2R2ALYP1XkGTLbovPR0
cZyyEobEPtMzXP1JTjJetJwhyX0H5gX7WHQeDYpDNsLIJ0RJd8XDMC0bnW3r9ROg
ljUcyQ7yNt4hYGON/vwcQNdOeBliYsna1RbdPzs4/earj4RPCZjggtzNKhPuLe4I
I6vxtvmcFom/J2BrAHufnQDpKIg0zp0C7oZrBKraKJlDeWSP1PE6EV0cmnlLhuQb
Za+dWNxbeDX/xFi2R6moddgy57hSFG41JUqVUJdPfhxT3mVcQoaRT8PcUW8nf5Fz
O9rVWOjjjupY8fcpIMcRjQKL5bRABZHlzjUlw2Yjo3Lc7GbmC6rUm094IKGQ2r5T
Wm+HSvHxJwHbIJ1/+haAJ3Z5FkHpDtkt+ek5Zy+weYSIzlzWmOx/OkhzfyLF37BI
Hep2CLOBUbTbXVosP7uMp6Eg4+Ck+MX3NeIHkVrrZR32554Cbgqm2CwkpmejrZ4j
Wyt/8CFe1JpmDHV4uqGhQhWl7B2BenwjiVE/2PKpCD6VinUUAVNMTLwPi0ViJMfp
92nNEF0DdMJBjeGhkZdwrQNIppN2/3WviZ10ir4YXjJUP8gDfjdJEKsc7HGZmBRz
D0q6fyDOagjwsFrxpsmpV4P0XuiVWzqxmFTk8IF57fz6jAvQluSf8p9FaZD3N+tm
FzuQU7m/w6VQ6YbIvY9VrMsmI95V16FZWmsrBRKRoly89wctqXKUmev/HuFwKTVd
p9rG4oKqPUT/JVS48hUS3GenyCu0X/jYDXAEFIIqwcLBWupim9UQ/O4DfwNy9sN7
C4XYjrGZ0ymiRWUsUn/N15wAtetE+gFqm46k7pt5MbEl/uLntNylEYxZH4u3vQUE
diwNRBIdzo7X2SBzc01TfFm2akUJ4B9yxj5OdbpKeH5asbpOmZCe/rEtEynAZbJC
eJ2gYqmP1p1/YwcsnpOUxodyi/CbsqZG3iLobCrJ/mtZTTSaCWgZO00U46/IeYfo
OFNqMi6jAWb/vKmL6vhERrHODg0lrlY4YTIH7HZgYHNTuMvOXDgTtXqPa0HNpDNF
4IW3brD72jNMV0BdM/kA9ufq7OBf9PW4ETxJKJMN3K3zNaWbWJqnYqildHjGYY2L
NLNts6ImP+tNlpoJbDxqGsXvRvWg+70VleOC72/cd6u279IwgKQ6/X8W+mc+AQfj
XL1FoOzxLG7vAM7x6hWODHYv56LM6DAwLsV+oqfBSTq4Va0SS8Eiu3B0krGRyBeN
G+F+bUdh1wAE+jdGPGEp9xcPCXvhzZOYznkXKmuUwYT+90Kr6tiEYJ+RLoXP451d
mTx5201kOp3ChRrXMHfe+yiQ7y0OjZ33/Q+f433GLTHTDsSWk6hGv+PlJvFikBjA
5HJr41GDGDsijZ8n7oHI/UAy55eA0+x/P+wqhrxAroda6LuHvIRoxv0sGEHtie97
ZfavxAYCZyMe7cLSqnWHmskWR04aZ4rfHPFzflwS4ndhvvaMUFjVKbT9Hf8dpcA8
37uFG8qRcsjgQSg5vfhcPZ8Wvy0OPYqs5IxMhbmj4aixJ0I2QSAxA+lEPytvqdJT
V9JL8c0zexCRBIQEnmuj8eh8KNlVfKY7eo4uh4046STFlrEHG2iEgA3Ss0Y36Xxk
vaqpwCdViQ665bNHFtb12P/CC+w3vZVo26rnVTbnRSg4U48GCtzDbJIWgrfIEKo9
1XFl8W4wdPcSXSUP1YwsKWqYWx3+VijgWovrJMdEBbPkLSmvwHYxGgsG0418AxtO
4/YNwslU1RpaDtq+hWo1HuPO+rsmrPuB9fil8HutPz6nYTb5btN7xrwSgCbOAelO
OFbWwOBoQCl3WknVmE0qLtOX0In2CQ/PhY/WlH8BG5hvaBIew9ICZ31wDW1073lN
xbwmb68w6l1GRir3XFu5JSpttWpIRw5FkJ1H6Ckc7aL6BsYFs+2laSepZVhkB8kQ
EAhHY/hSd5ICpRM4ux4dKQ+ypYU1vVv/bdkDGQnnAuVwe2fzXwE7yOIj7tOnXcEW
A9b4ZCunoTCtBw0JYw8kkRjIplsuYFeryhAKHxjbtALr26wUMLbfYa/Tof39cxR3
TLmaSfBG0XDHjWVql2kzH/MNqN/i4fXdLkMJTKQZ3ePGUZY4j/y9ICOYR7PG1mcj
GGaEhW0f+cIjH26EeKw8iDxqZHd0Vz9H/hUKxK16rKABltqWEmQA1leef8YkC7M4
LnOR9kkXB0eYXNyCBz4Wykr88Ed2WBRwDbij9OOY0f75mUAx+vVKcUf8C1z3V3qf
rC3DxUHgQF+2++rTDmS/qi5pzBNDf0UfFkTxUlBI/bHFiX0twtkkbWrvNV5ss6UM
vKwq/VGzDmf0LuBwXu3htVIFHlceco8UhLUVkZnjy8qcIEcfa4rx6V5g//yU097o
qk8XNn2hFnWqikIG7WP6DxkRW48kNOPNrqCoITICDGmyi90H1W5D3+MBjY3Ec1vZ
4Y+GXlbVoI5fd9lXiVJ88iNXWL2xn9RF4uuLGcdWiKahV+WkRaGL34/ly7tifsn5
cKc5cbm0JY9DPXW6h5ALXHZOnZF2ymnHEUXkM2MmrjA4UPDmgrcP253hXTQraoma
y4a7oXeVQRuS9ATYS1mvZ9IdML4nG7ab4i83vaDWxppri3q9YmKehpgaFz06yDk5
okWSS6comXipmFwA2dzZuTFf4/zVnLcQ8Ji8phMyJB9a2M9dAsmTWhbhI8BYwbhT
ME6C4Ti1vRuXXibEjHztgZLxhG9NippIysyYFkTvDbQl3DKU4nRRsOoBYRD9lcHn
lKGaJ4gBCXZTYJn8pGul+uavCqRUWMiYrqp/Im+KoKKW23U+vJORk9A+BDQ71Pzs
mumqTQX2656lxEN0WjclwfD91RGy+TndIo76tNR6xXQWQsmHV50XaZ4vWVZ6TJNo
f6xdZVUeJg3Il7HkpGikm6Y9tYBj+yexFsn+1i0beR77q4DRmoVgxxJq2qHbfGbZ
++yGVXxNFlqzAvOYwtUeRm8Spf8JJeYG/QkUcXdnyQRLs6sccosKJ9D7/c2DmsR4
8q6d2OsxJEvAXkbHUC5fwmltzoIInlJQHxhjPIpvFz6NYBevzFH897jMwfjprh9t
46ni5GxUov1B/lm2JPZkMRbWhYHQ/b1ozRAU6AQPUXWNDO5AHED4GFGetJwFPaNQ
piXj3SaWlFYbFAL6gIyI56TG4NOYI1pKJ/edC2snJnAMEv1KxcAOeZ4HpiSpi9Gj
lhf3OXLCJ7xP3IGFyni6Nxt408FeuTqv3ejU02ir6vrelZBap7hHS2RtfLqeUCxh
aaAzGrTaNEgVSDeyplh6HAsVJNQBJXTsj5MWDzd20/A+x19GxeMhft9/pn4YThVI
tRSBaHCT3ZTQ/oCjbeZunczN05XK6qRuXLM0+R59vXQCB0lz35nziN2n7lQCfdi2
CUbN7o1Si6H3Dww8I+i/EK59cmknTtDGcnYJ4fjT3Ih/6VkXjKTcWmmZt8VM8VVf
Ok7ebqKA5YTe1hOQViDWdINU9bJltLjevU8PndFkVtilXcFFHrofOXXyfl6DSWIn
ROptcjpXQCAylaThTyN0PGGf0ZbqW2cJgoHGWpgFTfFmBMvCgHW9EXzte+KxmPAH
i55d1NpXRbqPZCKCJ+TbpoYLXlhwnMWo/SXDY3yNlAvhdVb9e56YFHYpZNfaXG7N
keU/S287ztQTHjlryp8qx6Q+KVLgOtGDOUMc+KA1QyocmdhD1EkLbssA9/MLXuL7
NpNYlCYYOqNRxg8e1okKoFerSPIsTfHoMGLiK5iC0M54+c/9ea9RMqe3JL5rRfnD
sLNkWdj/+imbi86G9tZhSsQj/UYnfLXsutw6SnaCaMHVbmrIM7se2TGF/DQej4PS
8Uwu5WjWtwECMljlxkEnvF04FnyEXe09rE+XBnBf0CIudQTaqzSQlgNgoFLzee9/
l6fWDNq7RANKQostrLnkEXucXF6epeQ8yLZ8ai4XaYuh2/GGDlCxmjJz7nAh7tUy
cDwVuO7igwgqhSQn74xUTl6dZ8bSGnkuCLkU4KQi2WUR1Id8smzgTQDfLL5vZf2e
A7O9RF2YfWwpKgiudgxYsZsnI++ife104N+hY8G0htc7GjY7cLOjQ4rRUmvvIYsu
+/NSGZi/73gDerbCE2PAx2aDz1ywXdwkJoHZCuOn3uwwMoIVgq9pmUq48geTMejF
0TteBHvb11gm38sTyYpClMsgLke9Zv5ercP7onvZved7tsmjElTt0HgyiJWQmJjk
VR85Ms0yDdAGSjVr5QV+sQX7SRoKwAj21YBqwKiozhmHzbiQXQfhONtPgvpQ1K3D
LAc3BD1AGY5BsHbhaN5MOgFtbdWfGrld73bTvBgxdNHPgBz4YZIlIbKG0QsTrUmt
pfCCVi7KC+6qE4GKIr0VXulKNGGvB3L6XpHE5Lo0LUbeFUiFcNc/yNiSXcc9dP3N
zCVoIPMKo8IZ9G1IVx6DPDx9xtzA3w0U2JttgLzYt6U=
`pragma protect end_protected
