// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:25:49 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V9oTGOZQhWxCH1l337H67zJ+mA1MtsoIRAeoOvjc8ABGASlC7FjqF1UfdqJ+iYHM
XoRwhKGrrV2gx2sFDq2q5zbMFpvK6+cyhxCV0VRtjrBwA6Ng3Tt/XCc2p3Xl5oV5
NdwaAaAjFIDW1CDtyypThHhq5JcWkZX1khNBXvUgl2g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9792)
Y/938i1tgxFvdCjgxorc8xc2iob5l4pm9XSGsrNifMTWfSGeAOFu4mNwlcH+yp0t
xr1gTicDa4+TAQj8AakhydD0qanDe3f7FspbExcom8qPL38I4SF9t4FsOCR7sDL5
cAlWI5Z3BNu+CX2fqUoOQrmTuGOY7slQDeVlLHVOsq1gD9pl6NRF9dlmN2p7Ubtv
gHo1ruzNATt9DfuEWk2wHBaAOKuYAmPWqVZLcamlwBvjONSZS4LINTeMZb/37VoB
7fb/KrGkp+Ts4pfz/FZ2WmoqaHv7U+MPKyDAJahfgzefFemhVgZzI9hQUw9kkYrm
twWp4jWYon1qoNVjXc8OjBHTPU4/TRjpbReYpHz+1Hk6zZsNSsnJYITQOrTZ2pHt
041Lvla57buEP5fYW18NxSWNQFbcfkS7l/y4noxs5TPCeiRHigiXpcSPz0fTcs1o
oiJW7MmzgY34WLQu3p1roj66dofDLwcgoLFClqeWzfvItnmzbcRmBaf4NfS3hvtc
p3UvxYub36/OVJqYIwAIvxUwAvH5Gj7XT7CpU29MSYsQBVn6PaUMw9ug3O7BtpBY
rqZ7CdQ7UpS3QquG7D//lS/yTF+xJUJR51ZPnYt30UnLzL7iM5c7HN/NXHQeOigp
PMLHPPThfHNUSQY3NVo9yz0b3bXNCzkmbiAp6Wp1Rj5XQJZ35BB1iSsKVGWnqN5g
78OfsJpBP9hF/CF3TahRbrIOP8Q9Fgw5SqNq1K5qpZODqA0qBdtGPqvBm2ijTW9W
B15qHYVjT4TqsaQN8NId6DdggR2q+LauzG/4KUxWZN1FgUggNEYzQQRVsNr9Mivw
TNPROMx+CeIh6BeUuC4/nm/Q0C/VWuEup6DUuTK5fxGovmoDZ2kD8e4w0bykjDPK
vJ9b1qgwLsjNXM6sD2UmDaGsfdw5CGW7z6A67BtQaWV3j/je+IboWxD44KvFUdEt
AAcZ37huO57O/aoXDS1yXFqr43S47hy55gQ9a6mKDXTK/MOKAt9hQU66b95hItpg
8PJ7UvSIkeiHWzp93NeFWMDIm4rELIBP+rk4rLX3cfZYNPpUEsi0r1bNNqaOAoBj
ZuCzn8CtQvJ56ZRgEmGDs+MA4EjX+/RqahLsZN8PVFkdR6o+4vkETSUyXwcA47cu
VVrJ/jQV2M9FZdHmK20JuumzGSLDlCUspW40shkw//YBqP0XD2FvVKaOz8wSwE2E
uXdVvanfyi2I8lSKwIh42vXbHrgU8CvNuNNdysfukgElUYlmQbt8fsSwQMzSk7Dx
1m6YPjNJQPUGaSk+gIjZEzKTm7oaVpQloucXbpuoHMwnL67U+gOnoCce0ubDGWQI
lqgGyS5D0CN2InMSlycySEPwOcRySb8q9tgQX9LhRWY9C3+YHDl29cXU7D2cWbCW
7KkZylC0tywtnRzXJ03k3v9q/Dzf3+QsFQLmQMhII0VTYmvehrztpCw0K89P2aQj
zX03QSLYXjOQ0GlyWnpwWT4808rxtXVddygbt3Yx1C+Ayj321Hz6tAwy21wl8hfY
zpF231gNM+18MUDeyvClL60gvMtD1oPa3rqi5nYADXQgaejiL46EBPOeB0ABVyYV
uNpnReEyWAYhNeTK78mPJoUFlT7oYxXpSCY63exYw3p6bAzd+4gRpyqDAfjFGK7w
r+tB4dCxbF2vL2DNb1q4JQXJTwrgB7hEsti+UW8YK6WwnoU7B7MM9XFNhzoCj7Gp
MWr27QlDHsxm8/TeeRuRB31NI4mm65saciowYmtbtwRoW2tM8eXxBYj//iSToD9J
YdzC4DvMw4/4Ps+JjQ0QfaKPfbcIjNXeOuU4APXcqH+d9oYEABMKrKtu0hGlT8eG
ZrDAgtY8r6S3nIAkxqZ5STs6w84cgvvPF36HWZ2GWDymqxl2RpUy0/wOkay/39YC
v+8+eRZ90PifjXy7q6FVi78rO+Kx5XkWUMJ1nvGqVvIn/dHR592ECYm7xOAKk0VP
Lm+sUWZYW9wwDO5OD9zUvUgL2g+O8+zjf/zUA/2TCBFowlFL1/CVc2msTzYzamtl
rXxiCp2nSZ77JPoVQECsDm21h62tMiUwfJV7V5AMnL9SK3hOlebDGoLe86JxyD9L
ZqTjEBSoy8G0Tjq5CTwtyK8wA+G6xf1Wu1319eTwqYbet7pAXk/DafF0sp6AIBK1
k/zfL5/cdV7ScSQXZmMen3oaydwdWdlCLOCCW4TqRyMsAM1xPNk6HvqVps3laISO
1HHT2TW7aj9ND0Odz/pEAL6N9kETrP6yhHx+Yjf3pxR1PQIpWMkofUu2yTCWhdGR
lzj+97X0eT+tds6fCJkoS5PaNHW8ey3+zsy+lvL705qwIv49e/thsuDvhLHIxEdW
SJ/gaSDsQN77Fro+p1V+v7haw+Z8gy/pV31VMnqsBJaeq7EQPmQl35+m7vDq/vj+
EO53Bc9l9q4Y/SKrZz/TilhG9KHIz3jQfxQYVBh1UmyqxwPFySQv1i07feK69nFF
PgWK2QjmLD0X33Q40MKhwXE4Bib+Li23nmjZsNfw7UFm1xkJcLS1XnYZAiH43VIg
v/Veb1P6UI333zG23Xe5EgwoQtZaK734iTcClqp5iwDecXc/LXrWygAMEUOHeKhy
8sWmC/SDjrZhNLI0PWXbGqRk7g6+WPbqFNeWOUE39TNqVm830Nau2+C1MMC8LF7h
eoXO+SBTSwHxmydib1d4Qau/sTMeKWqwq5irZ2p8+5H+pDoYcMYid/AitZQcIUJ5
NzLLRgym/5+KpY1AauLWQfkLj0PsGp1uqCY5S0YPKTUsZYO3TbG6ZLgMaU5HM8Pw
vtDYQ8wtOvw0mK5Xpn3Qt8YHt2rH86rhp9tLEtzHnk2L6hP7fUN6xAv1RnyBT0Tc
fihcBS9nmamzfi6qj3F5HCr+qwWofVja8xw9zTmWVXZUdsaUb/pshlezw9ONYdHQ
4DFLLQ8f2eTBc0M4C+Ip5rQ3UcHV0q3uP9fvU3/PIaiK7jY//S7Wl0ZKjMVqLxaG
xYBs8jVKDJeDcq08GzyLoRjCVFWLJaBB4Rv71Ez1BFh5Zi7wMpLIQoSJHIhjfoUS
dLxqEi8P00uFL/Aj7LKVePZgq3W9mBrzac3v3JgU9LBLzfudgEd5Z18c32yk9oW6
3KExEOuFu1Zlwt6Hv3Xj1AaYw6HrhT9K80U1BqGFB9QiWnZXnTGw3MbUaLVlBNH0
/7lJESDCB4DfCHId8Vwy5r4ROYaGZek8p1vWm0Zl9X+7gOmrbPnLmUGpxOJTvG4A
Y9EgT0SCo6AlByZfJLE3/GclIyD6+AkA5/wzQgZk5JaDjG0LvpxQFWg7E/k3YkZT
VpqBqnk+TuH26uZJVXZ33ttXnZt6Z+E1QyXHc6eadFJANR87ng947h227ZKDzmR3
cUECP4hE5T8LSJBhR+XJw798zACetor9Pt/beMxaPuvPmeZyhT1dbb1DAWa4mKhX
8Afi7SkgVwpSSIDULPCwM9CBJcvYLG9Wl6VO+sUPeOQhjnay4ddCU/+4uX3/hF5q
QrKP3kFFBUJs680yaDXLsGn/xMkaTHfHh3NFgZeCbH/niMhy3E2NehyoQ3qckc91
1jPrINHo6oRwOEb05AaMlve1oZhPRKTVoxsjz/inL9qbL6eZG2oOVih/+VtHQUHi
7SJY1AyC8J2ixfkaEMJ39Qvz4yuFnkpMt7qv3IYF61SLii6cAoT+VcqRtD76+Fuz
YwvkRPp4lGWWXVcfmJ1kG198270xeHNZ+v7DfvDyVoz8t5HkdLCKGJ/E5f5Y8kfJ
TCh9fUFFRz5y0sPun0IWP6SxerNIIcowSmxFkSR3l9hsDG0Yc1nWtcR/eKp4IhO1
ap0y0RIh8vv0TacnV/kETDYYy7+1NzN3fM7tNb6bU6fqkRLE3ruSryM1Hu/hs8sw
V44LfNtr0drLcBsaGr2iqXyPSDch2+EdA/abceLaWe24AyrqBTRHvP4pKUChK/mf
QSSR3wmn+4zCg9+OwbKfYhb6VdifU3fzlwsmutjdoSs/IVNex3F6NIDF4uNXnEm5
6r/w81OIhUsilKiYuBi3yTwjkGjQuJEje/mdOANY/UKiCN5juTwcHKi5HEAIaj5A
epcB8h9C9HVijj1uTbmN2ZkvJ1NGsw2NOOvS42ZH1Az8ouWn+LQQEu9YoEY3I3z3
mIbcui56tAjYooCwo4zvnWwq7lMf8VM7/JF88sM4S1jtsvETg+vXoRQRq/TI+saT
sUiuXtaRNstmEWP+rh8YH1dT+sVXUSNAwpEc4iM+0T6fe7Wy1jx4a4KlklOBhsnm
ldnWMX77w4DBQ8wBeDQ52fO4qjJ7CHXr2WYZOT4fqME8eAtPyrOV0sNUuJpqT2iP
jL3YZNIYrf0oVe+8Ixt9KWF02U/Mswe9I1tFNf7xAcyToM6R5gsAve6FIxd+S7VM
jcN/I1hxbMC2yG9VzuU9cIgldB049Tigx60S1li0UJPA8eOJNMze/oLE1nSps4l1
BYjTsq1JKjJ2SWs7Bw1M3f5MpH9KlWF7PzRg9sQQLMUtGdn07Ghdc0ljNTRVf2pI
0Ru0chiafw86bJm6vkISldwsKvCP0pVxjNZ2OVzVya4in/DZILpzHeLtBYZ2LaLl
n328p8U/L5gW0IMrqQnoG2DK9xJJIelMzkmgtYPZjgopEUkoKw/NYy6ZdBvyM5Oz
5HALCREckJOZWxsiX5eFSMQzFKr0jW72rvT2h+QsyXsAZyEKExtZ06CFe4lniQ+4
6jQcepTLDuUCUVwON9BYOrPtynZ/gWe8/DNe5kcrF15aVVsgMqivcWxJcKM+d/uC
tSoGtjcf+t0dWlHKzOkxXGCRVr1r1hkw4tjSCcG7N+/UWX6SiMy2kibvhCrmyYC2
taYh0earA2TvxrluglWZeiHy5IUKfMaKQn4ajT/16JX0Sp46WHuyFqApkoTIV/7C
CLrmKpIdn1Tqo6hcqDV3Q8OUZObqtxPWkB4I8rb7ED/OdPEgjC9okxpob13m6zz/
JV2A5nELM8HeziKgHmuQHmNV0AuSutNu3J5Zaexgt/49jlV7/fJ38F27NKOzGDYY
LEpH8yc1pWy5tR73TQ+JR7ifnIr+09PWBFTzK2qG+3TMJBZRvr4z0lFK7lwyVZPN
6lZCRTo4RptTUYl3xwj4YTQeZrFGpq1dsSEqvOURsxlxMEWzkZPPw4Zuq1m3MlWx
hVn+vITI//3/6J7XHmD2nAOl3SajlNr+MfVkYbyoY5cox9exu+ZQhubEV6T1KU/Q
AcqLprlrgPfw5CCSPvXrG33cCiZT6gLqtIaaBO/dPsrnSvhvRFTFy02LH/55C9uk
R3tMmit7TsHk1eGshXXz7I8mF0GqnkhrLtNZWqPBG7FqjMFYd49gEuM0ksmvYXag
+oUWElLEMVGqbx87n8qjVU3whcmKen2xoMhThBsIXDBfC5h770naFu89D7hUGthk
r+u5yFBMg83N005ydEVrnKrETK8n2M1L+dSJD9V/Bggvy1e80SIi0Rnewx7MPEZc
9kS+nMe8gkA0Ug4xsejujMJ0+oUYtNG4VEkWeXpnfxxDmeacws+WOVPuAdJRX3x+
L1SyVIY0AfKyVv9kQ0/ZdDgqV7J05+1B5uUNbkT3eGN6/xFk/OYCu2tpbwgaRB9J
cs3oAAkkRW0dq0mMDu8laocCYSDAuoF70y7+HvgChM5d2NFepkbn7CZ6vl6SEpOK
NkRZ2QeLZsk65oJEbL5x4Tc6SjCZvhT/fl3rSbAGXC04wcFa/ybyYLBoK1siJNpy
Fitk6ilQXjyGhRBC1ASUXtDrMKtsoI5Tss4tnIQuDnH18P6909FYEu7uNOawdgyi
6tiN6BFMa5ruK1Z33EHgZsmdiJtdnlccduaebQJ4NXRtBB6IsprIQTh1Ha2xz5QV
FuvKQZPFudyw/Uu3aHrtU3DTJehEKjyVObKb4IlV0matGYKC8kP/JR3Y1q9fifqh
aGTma5ANZPiNx0oYqLIjfopOx8F3QpRiFiNJwxKnpPfapJs1jC//A1wVcMqSMV0s
I6qjTMgt6epzogk5zymbxbS+ul/C+5rH45lNMCTpna1nwS1tOpz18SgO5KtcMEwO
IUEL/VmqIvqQVVei6EWtlVAwG6mpcOfY+T8xah9b/Hg0KdU76XUajU6FbPTGugKn
b5cQHXzzKSIzFRDVUaPz0As4bfPUDd7MI0pT1X/zw8WsYK98oNY59Ike6zt8xwBv
gttJRhZ3hBZLXOt96D11+eWKF2DMmbKX2xqhsmLARcwUGhOkUpauou+ma9GtnznD
qRmQEu5U0rqj3Yr+ccmXPvKPzHeMOr8mLoiSE9E5BhUD8SPuB+cqTHw0uTj6Y8yC
7Cmz15UhdpShY/rMUoyCWPtZWBO22KSLZ2CC0K4G6A2Rublaa6fbeO2r93wUhbGp
gmV86Y+DNpJ1Nv0VSqc/deYksaONRLJXbWVUy7ce+gb9JsDkojMVKb4RBtfWhifi
asM5Qn1ThsQRdZ4f9MBuBkubnFz7mERjfYzwap69PFAj8M8b8BWXUI/2+pEojvV+
YVAUICbBUAlcAiZQ7MRrOHSlAG/lEFKOQiygyHCAMJ7F9AmdfeC/kcws0zFLiJ1e
yg5SeCvXYIddzViQT5zeWIVWnFI8tokXX39/PbdQXkGzTkSasQm8tPDZK/lW6Yau
GOme2pWXdRIqHMY/jJQk8W8gFi1euZz+RyCa0/TrWfr+59E8QjIHHBRXF7dCxYcx
JSqRgiFFMVJX4T8QEaFnF4asktxW/lkeqN6QlkspmsFUeqClj9sR9rSNQIP+ze+T
K9VcEsJN+XkeDokNwisVuxb6Mi5x5TCQCGtUQtHnCfQEpkw1Z99+6FX372C4+Cif
WRqHFWM2K4oNmtgIAqAdDerRuSFOXxKsv2+3hDv4Ziu0ugbW9uiurn5jjXCHYMGt
e72lr9xMNGY/AnngO2BE5mUDGY/XmCxMVtiXFAE9GX0oQqq7Xzunh8/tpjilavEe
IMt6M151h49Mxl8Zr3+JfjYZ0uYH5bHOTPyw4O6QOo9R4XJkXbVtDwiO7NG3US9u
DWPIrCRosid+Tab8fgU1y2E0fKDOVvxUCYeSEj8BDIXcoD+Q2IIhdUn2/f71gzSJ
eS1SUvIDFpJ7RFSlLkOzXzY7Ftgt5WOHxY2Kue2CZxGv3YjAFaPXwUtUsoVbUL77
RXZmmlkKZFL2CazJpXB0tOnhaiJkxy+KldHxLupoTkSI4twxT2l5DwfF/3gyvlUi
JGXeRcLkNUAL5zYZx+G3yiIVEtZhaQRyHxj+ULsmD0rd+HDV3haEjltkIxQJOyJE
R01b9xMQ9Tvkd7jsy5oJXwdi3tVMwo1VJp69q9NeLfpyh0YPz4+lXQQ2ODJpNACY
iQZr71vZ2OBsD2ijkPtBnmhjPEch5V0K1CrAsxcEgXx2ocKuCmUK708dBxDrQ8Yp
MI4/sRXfYcH5BBOhNDA2aboBvVNu4lZCTQHkjmw9JWb6A536i/EZz4MZf1IRCfHu
SVFu/T+bphhjSbcGl5bnilEdIUaj6a5bVR13WFMGDVB2iRnTlw7Dg3WZNEJkRwHb
P0UggV4RfsVySXVLwP9c9zoQBmjCkQ8eEp1UGk39Vxo51OebBKnsnInJAXFeGYUD
NIgd3PRcDn0GJtUPYPcLESWXrE2T45gYgq5GRq9wVK/U5oNU2Et+li5R2eCvr0tt
2mWXkqRPkbyRn9yHVnUKsDVK79Cfezp7gJY8EZwF4RMglAoMIj11+U67HjeiBew0
x1rwC4W8UKs4D7idpO+i0I/PPHP2AKSjGwuVbKikO5eIMKiLqNVBvseZ9vUy5Un+
ezyZYHAVJuFns7fbmodkB4ry8p1UuYL1x7vpY1O35aWIBNz1UbiJZK2UTvOscrOX
ackMjRCf3sWdmlYMtlBTpfsrJBhQeqoZ7STpIovpqpZV6EPbKCta8IE6xZbsNxtP
gaHUgVlrYXPplm1Yj251UkH49TbGsse4gbEMyBgHTd9Zt0MhJPjzETguVhiIKBtG
ualNtrfTB5BmEwOEN0TR+RwM/ZeLm2kgJQnhV4XzCfCRLeE9TbuwfTyChsj8NEXP
SBH8UkYyFENNd6uqEnARqdxGIXKAyptHXjr/C5jE+u0eCcl9ki4ldtlIwkpUqGJu
Fvr4NjW58tilikQa3oYykdmfxZTDlBvLZEspPHvNba0c9McENk6u4Y5HySf1O7Um
5IhvSbusXYVtY4yXKjJuuAMoLX2G14LjB7F7kG0hrU/sVNDfvBc/f+ioAx7Q775l
fPp9ldHksZxJWELmKYwCEKPA6MClVzJReF71Ryp46kb+kuUjHNfEsFj88tx1G8nR
D8zjDVwnOiBCQN9rEQKgVDuq/X5BjiW13NWyRvFw5iFZTK+FKljfSaIymE443Ekc
jzxAVZtNFxu2gmoZ4CtkaLn97kWZoNCechPbZL8PbvSRvHocJ9inb2d7j7XI/kft
xbC+e3+BfR9psyqYL0Jy8TlHjPVXXlKl5b28pgPUR2ILbYUieO7PHDwQheBStnCg
32QVMO0gcUG4rZsEGLZTMBVAJsLaUVr/r4caW8flVoskuom4c2Uyv6Qds/Kv/y32
qui+uJP5Y3t4FbVWiR8bBP7XCcK06SkubFnp0t4X07EQMjbuijOAW+OdVTekEeUF
u2K/OVUQbt+Ezxvim0idhgPbMjT6JjJxHNXYZiQjjGwAuNM+1TLqsuAjjHENie8I
OLxN0ePCePPuBiiIcjcK6RUDcflKrxQ/rXtBOVn6vIuK1vY0V3CmcwQg9lqOWdv7
8watc90jWMlvhQhJ2mJc0Yk2Mnj7jSpcFSwPO6VBpd8qi94tYVzXwEYMjknV0l18
3ul2oy2vKobIo1N+XdXOm+4ioTgvTxUdsJ8tJHEJ1PzokDHTqfScE0ckIi5Pczb0
28vhry7iKD+Ym++AdHGu5pfTC1g4FRW/6cXKp9/OziZJJ7ej83hoE+db1/MrU3lb
V4uYDDQEQ5y8aSK3VGcIsM3gZPN6o9xFJLfAoSoqh3sZ0zumG4rOtA6k6cBLxoDa
VC4qs1LHoV3L77LIVv4d5n4jfNJJ/yM7e5Dlclcy/IPz1/gKs/f/3r711XieQOrT
NHqckulo6IVONU0o4DT+Bi7r9c3Iqlem9MY2ANuC85/EB/Zbgc8jfM0hcuebCGhP
5cVPJBm7eWwv83L9+bR/l6JGpLwgWTD8pl7a+ctsK5k0y2T6nYbfk6cVxzjRch/Y
VqmoMBN15qvBTC5a1vMJdup8iinu10HxhqoW5swVz1yBO7366yMieKBU5aZEu/PQ
u/H5D22yWUkWuueWfwU1yNwtXDRwwe59hp48+X1bHawpHoBd8TXc+hZKYqMN+HVp
63PnFFkgIudcBOm45+le303Gm24tM0bXu0U8bKMJomBcyCJjX6FF7PrwTfn1LOYs
pbescWV0Xpt28cHz3CJwkAgs06z/yEr/lq3qp7Bcx/C17MtkpcD/4tPltkhg4v+H
WA/9RCV19n9VkFO3WKmQ4va2N06RrkUwvNQminbHfvDfJeL1IUR9xZIG2rXhT7g+
oacAqNMCC8ZJhyhpOsssgs8m21/EL3QO/BCxA3uJuXABos/bKlbj9Ipj4IP8Zwdm
W9nW8jL5CIIav3sabAKIGCWyDpzV+p81BZ7YpDgR6G4tasBC5TOPU8RdKZH0LARa
psI4cMF53dPP7KCGuJPpoCYovJxqw9UtIooBxKzwWUuorStvHX+2vG2Eub34EJNf
aqsE7nTiHHA44z9H48gnffsS/blnAwzqH0wHztT/F0HT+04q6tJ66D/psfaZvK5h
TBhJrQeoO88RImPk/fnVEgJjS4aa+6xnuc6+lvBGTbyQW6ogyn/ANBkBLOjpVVaW
CR16LCF/NP5uUgryWUJ3cQbFnXV6BMFGg/j44WmUKNiuEHp0s1EDr7LCDWJi9ROa
dJlF++dwwy8/6TR3zK1qxeZ/nIwAyrgRXNtRZffRh9TIUIBEnYaVJrqJgFXoV/Yc
SzSlX+XVH+YhcGu/r1qQnmokR2mDE7ytQOqOkfSfdJpP43jbHqPz45BPwYk+RiK6
1eKxLZ+QAVBbZGRUCyR8fSRPBEgh8kI5oKBhkMEHFALT40nWtWHQlEDU2fmMrs6N
sLUj+4d75jWGU09l4GNoH/D51t9eQZaPewwmmeAvLBjHkk43mOv9N9iqZU9P724W
Gw62H55g15UnqRZpOgDM8yssgHEKwSXeFr9C3SMTDDF//tAsGXLp5s/i7dHn3hL0
NTmqADPDL/zm+8Q9rgBuyYScE9EuXaxy2gcwD20SwQY8yiVYqQypFx792bottevN
geXXiN7186a/EkrfJePpd0gA+O74y7v/vbiksXbiCmhZKm9HieVGuqF61mDEUGwP
bvksUViAu0eHYk4ozJnpKqQBX6Dmy6AbDK6qW1EPhX42+9ZIQesmpdRqodl6XYfd
i1t+DfNdox6N6wSuBCVT+icHAb1EeEIjHXwrjE8WGS8NNarFw4X394zgsIZz/Iz1
HoREYbhRc0kEmEF/Cbvt4el+h1aiP/0P84ala+MsDSAGlpTN1fNAaF2ShgH3ZgMz
yfIVPP/S1gIB3I+FHqEgJoQ2QWoFOjrNMfRNYToL2mS8UE9Am6OpdtvNQJibOWFS
Mj7i97TUoTeHhXrzNf6tzMYny4z5oThYpaeECptxeK2xTWL681CDrx1jMeDx1xm/
EdqFgGK7gIR4fdDX/S3e4ZDYdSQIzVGuyrlq10CqHLuTpos3L/6Dqq0D7AZXPtJY
RtbhGUrQsOsKGJvn+VzhhW1guvqxAPixMLFeo1Felj5CFzkmDRdqDi5b3IIHWol6
oe1iBsN/tYPqH3MJzt1MaH4O1NMNkobmqJiE5Sjapw9lgi3dZmWJLgYjKuR+8BNH
wExMEC3Ex2qa0OdrHozLd08Sb0OCaatMov30OyRzHdE1iCnBmTPeIbmtn64kxO25
TDL8OXz/o8j/nhHd97EJEPa1k/X+zF6YmKg7hjfgeId1IL6zayqbhT7CaeeCPMh9
xexVb1YnQ4bqqPzFi+g5ZXFdgSBD9zBpSLbXZaqNfi28B4ZYLBZLNfATOyHETy5k
owkjoIzoWavjPywx9G71C3OhW1RY8dtOvmbs1GDn6bFRv6ZeoeueW4m3ISZeY/gh
SODDG+CkmyRqZeJ7fyAnpgpcwmVdu2IOCZdGix0xFhsf3PrJlQDrQgVgCP8lqXB8
mOJ4InQmtJhqRgPQ3kf2ArvA4Q8ncwictVUYh7+UxrwrXMaQrWk3Ln8nJC4xm4kX
ZRFCejqnTLPo5jmut6Cd/eIgzaR/IodAPj9RH5/4ki6YYg1v8hl5O0H9zsq+G12m
Z6oBTAFQPPapyifDBhGKKyuGmBLhLeXkaJNmin8ts3F0SicgMeeCeV0XvFihsQ5m
oKnQQoeZ1HKxNEnfRjeA5uIMk1EMDUEQMbCmJenl8L0sYUf8mpihpNosozt8Oamd
jXm3HHbSDu+xhIZ952Tl8GsyWmDmkjh1AT4npdAVppjEbPsGoR8SE1YxrvRrYmvi
b/JhfgHA8AasctaSoEw+HQbkO9fbLJyI1+gL8L7PWLpM8UGBPYo6DNCGjXrzUSm1
zscufXTW9knBvT4iVKQYJC7i+yPOfjoRYhK/eRG9pMNFttV4KXQ0MRlDlw/bNRYz
FgeMZ5vF1xepnKZe1KnwArmnSp6uPmu1rygI81xZwAn9r0RrBwsD2emMxNvN+IJM
/k/hUjSIXoJegb6wp4dj7P/UhBXCkMP1v33RHH6WqXBZSWQ5E7YQmOOxbWQJVw2W
0W79TO0rzxJ4fJiSB4qL0pRkcoLqlogd+JIOHXTay5N6iKew9F7C9qTfKxVM/8+E
q0yqJ27ZJYjTM8WpnZPwkoOqj99e1rH2Sy225AzDl3q3e0g51gSPMSR0esiay+jI
wlMGYoO1vcKy1UqybT0vhrC41W8s4sXir1fmSnYLDuFcQ5mbxF8wnOwVvfrCi0pA
HpbrrJvFIHeuIjHfrtqF3vgoLpv1v8aS/NpzLRxvEGVYRLQ4e+ayqQ66kPoUEBxb
m27ip0kdJlVJ4lk4Ls2F7R6YEJ/+8Av31AZn9FkxYVxm8G9/N+hukBxe2pGw4IEC
5+NE5HpFFq+gQbRKpiIdOzXBQu4gavR7azN3XB7O2UCW7fVUODH64y4p2FwEMDiH
quhDDywzOIaVQ35rCUO9DFLkESCx9IvFajXjfnP2iUrxRfPNt6crNRA78mQgl/im
61KEaS20oN546jx9DvUKuADZEMl+8GRczcYcHoxkM1BoJSGdH667B06U4bBaYBXu
3WYBOWXX5yDUbnbAhfH4ZAHpnUIkzHq5u0UKEKnFGAtdp5oPW9tqw0xD0HEY9zfk
RCkYTsTuaQbbpuqNKZV3wjhtBqfAHLOUquBVhj/JVvxLzpwT9yVOWT0n3EYH9xAn
mzTXAuFCJsCf4VDpbMnL04mvke0h/TsmfdMAPZBIZr55JWQQEELspKeT85TqwSGJ
Y+hXTzaAL/H6JNLFRG9zNiZmAfXrdh9eVqElpA1DjnqStb+D7TfvKS/l58R3c8X/
0Dtctahlw9Uho5LlqBKlrN0KA+exsxSH18albuIqxSd9BufrLZjkobRWI4gvmfAC
RllNXeStj1NhuZblKMWqPNHMsKEw7uexQ9Xl5oxB2MLFWdILsoYOScc54zOlT4Hs
1uO17p5MsPbI+wsPf1SbW/1/GlIxJZ4jCUaAU5pHxjq9EhQdYMvUz/Or7xOKm3w2
IEkSv6LkOxra/geFwHU0EgS79qrgPK9ZPo2e9AwesNIYxCHxg7n9FXgArnuzHMjt
Ky/UFZu3hpOEKzSAdK0VsELCBZAkLmRkCZx0uDRK2VH3Ydj96k2NwoKOGIp7l80D
5p0XvLBt5fAQbVtgC2fz1+fmghsottqdxGgkiLTMYRysnre6A2LwqksAEWWr5A0I
Oo9uRiQM0xM40RdxRKJtRKj4+kVWTQ/WjpSv/pouhj/sWKL0iL7+NSaJ2Ns5y4W8
EankA3pmTdOyGIp++nYTMZXzoCdXc4BYXB/uTSIPu3SZQFwUTfSruExaVx8qIH13
`pragma protect end_protected
