// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
YbaIJGdZYXnK3xUbWUn215piw6liZeLuOsYfAwPnqroxKZHWOUyfeBpg2WWWbL2UfY/aO9smiVEd
6k5ui0CD0Y/TS1Bo5mgR3g6dWS+0vWH6P/Logc+qZPJ4hsnPa6a4q7Y8McTkdTQ/Dzo4NtLDkQNa
vFey2tA8rZRHkEUG11ZJnOJkUJ3UhfzWdj+IxntBcdXcaRisYiQIs7LpclBY8Gdcyo/XFA9ypAwQ
q1HcIWIJsTqerZx9PONMoxSnePT0GK4l5E0wrou+h1uAk1l5nT4JYHS233qrVzkqtNknOKa2rPu6
6w4m/56E8Qr9pAWEdsmGL/8H4wNV0bnTFZHYeg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9712)
1u9NAxC2Nu+4tmqEqBh848PKS8IcixY79p42ORp8BJG7TDHdQkV1c5beYfSykhlvnz5deJ+bIste
HuaFqUM7oWZbIg0EhvNMtrrH8gOkH7AXYabh3RFu/pK30Abq2r/fLx/USF+PdO88nhiT9liuhleK
mJ2hTTTZw8hW6BLUZsttaQ1sbzv/mQMc9LQtaIPmYskzh472DMgUlD3qhqeAAwOFubfaoLJJIsiQ
PhbbbPDFIYacU4H1A26MnHdAf3hFASyc2eXLFAhZSo3ndPhAzWzH4epOl3DyjtZH5YiLHJlylCxE
ivxCHAiU1ae5Nuk1FuQ9HGx6C3HTLqcTQt4BHiuLvuGgapHjTRAKGXpEWSfSrrQe4UTZbDbU7mUq
U8MvLkYEG3aT1ugCXVE2Ko1Dtbem5eFQh799GHmOylRgaimIlgSC0NhtU+1ZxFG2ul4+vtC7JWJE
VbGg7fnZP2ty7Z49f3GZSqkXPzruajUV8YBglaol81BEZAGqxxt+X3h4hVESUrrUQlmXu7WXi3pe
IJb7d1FftA+VdRednX/q24wByJLj8F1gUgNuY9rvG2r0l4bLHA975SEXhUZjZmaanKUvHxc6GlxA
yarvWEDf29TnyE0hticHoO1zq/OaavvfRRd127i6ORjgNNHn6x2OW118UK/3DdPJCfAdEcoU7tVy
VaZ9VO6S+A4QljThUcc/PNnz3a9OI+bnf5pu6nQZO1QezZ4/Go+B2m0iYHiInIgb9bmMUuSgo3ng
Vz1+FCpdWd3xNCl+FAy4budYTxbdfc/phCZXHO3X71Iflg2oTGMnMA1UUIeuE4LR5Egmluw9CRAS
QfwO+9EADhAUur/D+aA5gHxhj4hXsR3E3E9+sXosTiHY5ra+fRlhF6yFgnZNJD7K5254roBN6rM4
VCfSvCkk4CJuxcySJT/cvW8i5u40THKCdJQn7Q+E6SVL5vgv6fSXmmsb2Hn4bQ7jg2BKbYZkpJtD
M7/4tF5PMTtHA1vrg10mz5KhI72k8t/II9WY/tFRf99ZwhshYeA+70lOM58cJWXweyjCL/enQrIA
kJQEZ2S8ms64BnmsDjYYLZXJwKTBclCFPcZoWWmee6cl3vLx+PM/WHLG1M4wQH8KCWpshYkC/GOY
jzyb0wrbSfkVWcdvRpQJoVvxEVT0iko68DeODFDxCI4DxlzLsKGJO3nR83SMluxVWio74jyZmBU4
0KVZdc0UAeJ5XKroHMPFSf1tUqW9ToJaEDewXWT+iQEg5bn3XPPJ50ircCnPZq0UR8WFCkL2ffLb
dSxJFnxV0Vdk/F0tneNRjOMF4V4SihT/O89w6o1swH6/AGa4QIngjRA6Lk1OJ2fSiea3Wk119s/W
5RLOXAm4sdc9lG96ik75Ym28fhFS19KjeS9YtqSeNNweOECCvl4FeUlnCSeGBFYTDBXD2H9rEqF2
zBWqCNL1jQhVWX660B+NC8Y5Q1K7iSdXmdo8NpXeph5rZ0Mrf1+WYT9a0hrnzRuxFK6KICVvNLwn
V87pKxGPnSMV0YVGaF1zqSmz3eBWGxcSdt1SBEYs6vU3pgz9mCTvofcroVXZ1LPN2YlErgOXP1fG
w5f6YsenNuprrnkqwZYlsYzqRNGvVugE6BAiErF1EgLT6SZ1ZP4Xn+bKjDFkygxn0oSlqap2Lin5
eKbZao8ncSgLsDOdS4B1DQQ4rgbpK5/DsgurDCJi0QZhBOoHX6MF2dlYMOnxa0xk5yzZ2hnBsQ13
p2u83Mu1c7TdRR+2vem4sDNIKgwcohqjCQPwe2+lX4g3nA3Y3bUC6Cq8HugfJYcgGJwxCpWy2n+c
XHMrzl3TlW/HRbiX6N5UfM5vYzxU/Jer16C/M5bHmbbcxwmVcwSA13EdQ+nNh6LGaCnIJde3ey2f
fV1hjHLEugl+vWYFU+d2UeXppvB36t+KTomRUnSsdC6qsjd+DMkPlGOuYFKJHoKhAzQNz+ohYBi+
kGipX60pR9p73tGAvkQ9lX5+fFfUns9CLncpuX6x+e7USbU/pjKrR5iSTqCRbdAkjVKQSN19TreD
qGw3Sc9KCtONSC4hH5wLx8JJ7bbpUPVGo/qETuxidtMghkeHad7jUUfAjguj7mGu5pVfece85T9C
2l2Z64b25qRy8e3xNlbzU14rPTZh1/2hrmpEOjZqdhlh1A97Fxi57FdHbbeEGqt2sUPUYXbcdPtR
0nwFeUQE6XwSq0CCKFIsvOURT7BsrXxPhUU612Hw5v0vTpz9TkSI4iA/wzj0K19MvGkpBxiVRQov
RLNplvYvzwWwWuj6AJ9P+8hCIFxXdBnOq9AT5bJiflJ7PHTC8Y97AZiUw9D8M9JHEYYjBeX7ihT2
L6HW31oahpXEIhEZKy2Pj8BZVea8Gz8nv3d7guzdhwJ/671AXHmShdXZY3hdUHN0GjHRgf3BZBUf
R5hRUAiW99QBZGzbqvAsLoNglf44B9x3IY2dmm4EwMNt2lxrFxER4TrIeNbxLNDStu0y8ASVLupq
SsBo2lL+O0iq0xy8Zt4fdAI6/MJ8CA0fokNkc0TsTI57B1kpC0rOlKf01Qp6iJLwguOCdLCexAu3
73d6Kl9/nv6h6gSAOAn5C1oCCUfoYdAJrNn8BtS9KjN09uNZ3D/6G/h2SiQQFX3rN46+Bq00byCE
z34MFWCpWTwHOYkfqatdeCHuR/SJ5KzWoKIu7NyNOLig08PlqLWgucCGseCpTMU5zaUUHCE1XIzm
QNmDJr4kJj+XyCiacftxmPD7z8TzOYDKCTEIh4OYeCXPKombQ6ReJees9KvFH36vgP3O9qZYdkST
jhGpmNKpllKCOfGXQSFjdxJY0hh8VWlpuZ/A1dd46FGj8rgQPFMz0AliyjlMfsigu4XzbZfR1KzQ
WQTZbLcsckBFqUpvhkJn9bLB8h9aK9JtdI2BnodZESiG9PFUXqvoeueuuCvCsQQGUAMiY/8WigRm
qgkI9+uRmjbFvA8M+fe8iytcfWFD/f2aUrGPHyooMb0oRs5dNKRV4UOwYHQV69Ol4UTRtVWKLGsG
4FM7pynzYGKlQmLn7Jvgx2wz8ftsZYcHva++LDCE2kznhrwpeAq5aVn+Plhw3XdfbIaRvs6dihoD
9gjl9SgmTyEa6KCi8q9JDgvNxe/kyk3y3NNbu+d7n496RdFZaYv/M5pIk8fVUFjYgLVzpuM8dRed
nPYMLgVoPX3FcygtRFNmcUon28/4gAormJ5qqWQC0Y16NxnyuU/oBYuThpU8UFG4ZC7b2n8f1zBl
Q7lxPMuG4rPLI3MnA2EQ4SxxD0MFFYb3OIIKjIywenO9STPhIYaVgqKZNiQp1iVQfF9hpZq3lf+I
Sf8vty7WcEoU9atHiAdC7HknVJupeCCMPOm7uLpAQrK1vX/KNREhRvbqzG6YvvEQttkyfgWv7swI
lIR4P7lgCUXjlNzXOoGVNw2IvIUfnHoRAy+hP1OyBcGPlRWlu9nfPw7O4M7Aq/U9p5njS7qnPOVX
wv+58xCxjDtk3bHqFM7Ve4Iqy5zW/WppjIH0GYySRZzRPxKgLOeJGmd+Ge7oMe9URESx3ouSDhEL
P2BqEm2Q7o1Lutw/Sk6TEsyMwSnFqKYB4LmC9mDYxycAeYAlak+ZWtr2vut3iy3/7DGtpq8EF+BB
DMlpZwMqap/+Um9pTbqYdiXEzRzM4oRfLzqE2LQf2GkxstHefJrAIzl7O0WVIBjH6QzAJHhPQZJC
2ONRFtocL7jQyh/sNkX3TZJHNJOTiqukAEYUfcq1rxfgJ+l01lhF8X/Ufaregqca2BNFIh9dPmOm
n/y4kzIy5qmTt+Oa27TBcIR8ymqaefLeLgJVPIQyU0ykPe+a9FAjrOKrCTTvWywYcbcI85atQ3v0
QTIKqT2Qxjk12NbTgltlaHD4VPLqSUBR6vmQ6fsZfyKZezunBjT1F0TI6K+JCLprrxwLy0tHP4Kf
YUOJxR8SS/kJ+Gvo2iugiCbh/bDUNGFHnihzFEfMH5Kg0mGdv+BuiSIKNypIvi8A3a20wnAGKzIU
81YYScN3JTmDJ3kAL+bpqZMW9Xj8ybxKQnB6iIiVFU//Hbqhqk4SPnuhtcEzhIn7oSDeKYovgQ/e
wCfutMWOuChsn/f9WdlDO5GAdCmHnPwMVWFyZyrkhgHZaU3YMZW3ag8n9Ey2Sd/ANPN0hWUgBnwg
2r7PO1yJ0pq7FQEXha8z5Yef6sfy3iDvzyQQ02NLpFIRofWFfawz0+4O/hJS0qSjVD4+Bx0DFoYW
Wkk281uTGh7QRJNMP4vXa4TP7zrLOcftWWMOEvXjEI7wfHEWZ6jrEjEFhOsEdSubBZeF+I80NenG
WpU6h3LP07A7Gcr1oaiZBAWA08jAruBBbQO+SOO5rRPWB4brBUp2nFU9YRmJm57fHBSzESolPmde
MYvOZ06TZ4I4R3ZlVdIdVMQ/Yl2ZwEOS9r8p2CSk846k1ZZRk1n/L8buSADT0DGr7/8fuLsCfA0d
HXcgpdlpBp3+/IdfrOxVL9w/14wH3cxFYWOIdRPC7XafppSPlRugpbcXQdWb90E/wmN1zb498TTx
Q32Fhb8wDAEdS1jvVVU9/WKLaqySotAXD0IBeitrdB7OJVhsh4P+YbnIBmRaQIP/K+2yBUrsIpxT
t8PsY9UMC9VVQPZ3Tvcre2HzaNk8wJfwKpG4910EIEf7LAx1AvcGNCezWikO3fKqFnke4d5dKbiw
yQMz+lcexpGtmRBOSa7i6sR56fR/1cMcNYPcQlAf183dTaoMctxvpA6/StROtEliMVaDubtlF5hQ
VBDuY0kns3W2nN2BpDXLJP91eRqhl1IWuC1LcP2lkJKnLTjVK1yszB690QafsCWUaylf7Kvssba9
n6wvaxiCE0wcHDZP8sBUguv4ExwzLcbAy8aRehJ8S3CSeoRq45iWZkzKZViL6tXiGKGU7pUI4PRc
r/TyFBGtQHMVdiQinokdTqUrJXFivZjk7a/QRxtF90ocIiD+kU6ciKvsKTXybp/SYHqJLmowmcCR
1ijSNmcEOOZzkZGUN8ve3CxCNHq4l8XA3P87NZ1rPgibUo9u0RpIExYjlXeavdNbe1B831jE9T0Z
CczoGxR0Gb0i1SvC4SULLBc10ByzbMb/5DSZlMGN4zs6XO5kIurwrnlRZhAiCDUWHOuvbuzHzOk+
xvYMU+R8RSR/rmJRsOW0jT+xfRjwaO6pZNeL8MPDS3+4eNjzZW66xRKrXGbw61zQc+rePwTMEo9y
YHoiS9sVghsK+IOHfCNPKrjBe9ewToDLwLqAeTlL9MHOwnt6eOC35iaCftS6oJMeuKp1+TFtBSV9
IoN3E2FOw3/xO7k9i9rFiWF8al5vOr8j6JJ2ZsTDzkYZdaew/Vy4jEzvPdXCZihHrMv6BecUzFIG
4bLzL6FIMCO0iv8ug09DbSpIcVTFpEgOS12iUmUqI65AQLqStTejyGB5TYN4sYw+xWjGLRWEgKQK
InSuqpV3lrAR7Q3hfKxR73HDCxpgkpbpx+E2x3wB6ZRdJ6HCO/A3S0xSFTns/PvDIVGEVc9JIzko
TQYiZrH1GK068ssc/I0tGLvwc/EDSj3x0Du7kfL0KcfpuBL0jYwxbBdWbN6Na2Q1FVJCLv9E6xJl
+LBA8wLry+kuLgI70DRgtEFGkXpWTDA4CwbdjwP/Tow/iVc5SPnFDs5xlGfk2Yj6KZxCLGGS3/lt
WGsrnGGjYkenJSsYMR+bdVQjmtlsvfQMhXudwkH6r2BQ/4BuLs5HqaAPVouc5Q8pnpeOL5Whnjmp
EIhPhacLLBe3pPr8mqry0013bpvIcP8s62QPYq7xySmb50bSfs9EeVlDvXqAnA1kVyTkgl/SsYU7
A5MPSR0ySFO0RJnG4Xhpds7Hq2gVNob4XbLs8sBI1ysgUl+xAbiTvLzvM3/IC1FTEX4Mwon3fegj
j/jFMCLK9Wu/7TMliygaU9gnlXjOVTN8Zkn1GhxPlXNDQaBt4YYbRlPTjRV2DR2+CW1ssSaYCSmf
KKgimw5U/tx/pn0U088SAA7Yx1R1/8U88JSGN9HUqLS5REiHx1iClAiDVAQy4i3dN73KBFNPNvP3
+CjD1PO4l/dAy0g0+/AZoWq6GRDhKPNcibBo7c7F7nonnsITFQ0jCKXWIXZbbp44IEKreSu1SNFj
8lIxM13paYGN+IiT1XifOFJSX8WFKP1gfF1voPvgF/wBTFyozZYyUbNoZv6K0hKwiTne+OR0la3F
IsmzsUiu6BmJ3LyhDkCBA+ENPgZS2nzC8TZAoUt+BuT2BsArVTio2ZWh5C1uPyyzcrU22guiF3Zu
RF9zoSUEl8tX8EqxxccIbyKLm/5DTbyEMp+ZnlKxc/neOkRtaFxpVyI5xhfdNOyL2Xxfmq5o1nJP
HoHtgEKr8UoJYMLXpdHU3iiX3xgNqPvbx7sLFWzWibpsv3aGnsrjJQjVNrdOl4kFbiZ3tkUhIs3a
ufUy4vXrzo/yqwLU+EhmcGLu6sPyj3NvuovY+gvwaIB4EDUx30Y5TldGSuzZjJwa6+NYhZL54Ga0
/sjGISinQTpTC+t8rZzXwcQrBaHsp0npcFfhFF+NCxi6JJVun37Oov9w7wpCiqCURKmQHDlNeHpp
EHpLyQ2AoRZYV4nh6c5jbvsZoYXfcpe5LEo8dg7txZKZxHVlyfWh1un0h3ly3KS6GPfGOZFeVyH1
npVfWNEKXHaB0FcKc2rJfcRjYNhL+AR/wT5sw/xdVkzibBThevZk/q2ypUYpkvIWwCk5W58KDP2o
41BV8tXpBTkmiqrux4Zp+oWxt9nNriF2TeptYeS5iS8SxSHyiDQr4i6l6AGqKiEkoQPwQw1q7O87
PSrN5SOaNwd5JLB0AyP9+w6Y51XjNWUoPr1f2fNiZFXUCMH6D4jDUFWmNvTyNLtQVxEPM6huyMI7
34qSVqpeE5bOeVNX5jTojof5OS3vGHSMCFgVYgBYQ92zRW7i2MnuTpKyUzAGPj1+X4h1wbPPIEBN
ZYLixwJvt04qFWBAEhWWUJU+bfN1EOlDJY/WOhEXp4xzf5ASYbR4iGXZkIFIq06eaPtRqG8+JjLG
JjqShvEO0Aoo+dbvd/lAVEK9O7+mI8l23TvVUIhSXXJM7JubGLvaYO0K820bKA90iayyYD980tdv
ydJsixkkakWIHkL3A/9hvq7RqW9ROGocAO5VtgsMztXRD/LrDlR8z2JDl0ZbsSIx8ZH2kriGC4Yb
UmqJ5th5nJ3IzqMuIWbb+0KL/zzpDbR94dwesNY8Ahlm6V90x5rKd6TIQtOw8wJwNLBAV0mLSqvm
kSmjXMzhehKtTD2u9P4VYgarfahfNAwiMdMX5Rv2s1xuZvCX+qH5Ms5XEpWqyxxK46AYcggzlrjx
5MRoMevbOynlOw6rWfK4QKCyjrnJ/CjlVksgm9o7KzA+aCDbbrOcoNtT70yGzmeozy3slUdU7lkE
glcmFlS4yrCc7pVph82PLhE0ADI/wqZ+dD1ZlTXCJEk08vnWcbmSVqnsOoGgKL2nSfyklfvfAvcF
DvfN/TxOvz+LTKIqXrNrGQg+AzQWkq+AC3aWv24wIeaTrx5TbyZNIiUM/CFE7jB7aI4AIv3gHGsL
oubqIYY+xU+j72dg6MkkT5MDHBybVrlDy9ASpH5AlzFcwV+R0F51TT0HwDSzSDtSpCjjK+sr2efS
Vv4bftMXz/uvZDfz33uN3ArHxO8MFqSaIsmTs9nntBAvrKlEiEek3y0fwDJ1SXCfsn2LuxIy5GLF
Z/YSEMIJDC5Hg7McvAn7w7t0kVdh9k1w8oDCBE5URlMSRfURDfVzPjlbO3TQT5d6mCx4CmXQNRcx
qm/j1tTPVz4yiZfLVKczTxXP/LN8Tp30DDhSgAOmNqG/nuXDirWgSR1S/eI1Uzldi+5pcvUabGtr
uHYE3hER6kBMr9KfV0ttFpVzS9Rf3E7WUOIZLc4HQaqpdGqqZpD2eA/PjFaZKt7xoKoKpZug0FxV
HmuKUGhuw/5DNQTsAC+65rUm7rXzJqXe96D+ZTOROx8zsZVYFRWad1f+QZ2WbRTYgfteq6oGNxZs
CuI5W9Kwka1swm8y4IgnA5gJxPEqWOTUm3/CfFCo/i2L/XNtRRePU/CR4QHYJIy0uj3RasilpdPz
9PGxEytTUEkAIXYptRRU+YBF0ZN8KPGUSFKdDrRv1mMMTe5OQQYyxHcT/1cbVrc6cbP83dq6JArj
jgOyNIRI1Z50KAUqIo6QdVJMJgw3IA+BXRY9fa5QqvRZIcn3qj7v5Te4JOn+xUJKn15tE2HJK5s5
5Vyks1BtgrMFuPh2kkhTsUupSWm7iWNYefWjfqTNYxGzlXR4+99PszYfXJBuKhwUC+FDILVOtVC2
CEcNGyydtQjgxFZTugXYxJ1SRXlbaO0uHaNx/kxoKpQDYDTcGmc3d7BrRhFu8L9MuM37XGpU5Fpn
UGKL+Fe2gdh0fjLdi5xkOVPa8wIJG9c+ssZiuQRcuuKt6P5ekbSJ9ebCGsm8XTX9bvvYZ1B0A8FB
a07EiwA2M/sU/CM0txZYYf1Pj97Vzha6PEb3v0mZVVlGkBLTnx9E/x561lgIe3uEHHm3uvILwHKA
CPgb3g1pu7U/1L7JZYtAn7gn9DK4Qh1KAG/1gSZxaAvC88aESU4QfDMI4sT30VANviRwzdVUsGin
OTXDqttnyxzMtCrOjiZZ6w3tKeYcC2A7yzZhFVxI4mTn0PWhvq4/AYGyCbHJ3XOYpVIbH0vXZatT
BQ9YNzX43vEvNHZ5BwjYSf5ODo97SFRSHlfsGcDEFwWahIgxy9jkx0SrUA3ApXS0xfrPDS9VZOJ0
Y/CqaWagjsSb/kEV4GSiBwda2XvgUA/0HCwzCGzkt+/kquZcCTD8EX1KF9L4DFWC98WE5qckS7Vi
tkzlF7e1uCP4VHVcZZ5xAMu96CBaMJqh/IKYSLQn+iCv7MJZ/o0zbBfDdyguakuDQecRndTabmGv
9Q68zjT1GUlcZGBT2hnOOPiwddnUBV2UR86+rla5Wis9662OaDC+OpULmOeiXt3APs4NWY2HN9r3
ZsXtBQVy9J4y+7zNRUCTga8kECyf3vLyjSXtEJTIqToyJ47aewFbH2duUjjimFz65FD+C426ySkY
+1pAexdEm6zr2bW3HAZCWM5JN+n1vvXdzJFi+oGjzRpy2rIalXIM/Muix5VMWasFWucCavCNGdDQ
z+LMRgiTHfMOPbAbwGrSocIF+mYw/f7EnrXQJZkUdRddWj65oeozhGrlCxby5u65OrhjjnCnaHBC
MYLO4/Qtnnzf3PFC9LtdZakApKCZS/35CqoOUYlIThjG8BhhY6TnIFwErsK2KJPmJ2Vw+NtWYwLY
mhW7V4vUWC/zqzSI/RBRjJ5QhOkYe1gH96sjDBZTPTnAwq2DylEd5mqM2cw41iR1yVB7yEPq08Pz
Enbl9N71xvfDchyg1YqRcMSxJ/7VqdFYvFa0M2shXC7dgjfeokb6iO2E6NJUYseXvcwHItJMrbY2
rCPyPg1T1VL5yyEAH0Iz2rGBNQ0xQDhLATirUJ7NydahTOX1415wHR68Lc/nZP+VoYzO/bblpn4s
XZGrsYSAWF8dTKH5pKozbbPc/WwtisZUlCV/HOrJPfKnVxKzhH9AYs68zqs8R4JTAMJpQKQz2xRp
K5PM5CNG7VEvvONXh59+cQQYhXEslBJPq4bIfzvgBJQs2qBmfs84be6VEAweEaPsD0c9jTUZQcec
+YkxJa/qCHkmLDil/DirM1/z+hR6mamNohmSVV8x3WEOb9tayb4rg4UA1DMLEBN+uGGEM3OIB7H7
UwIRycCpgj1kmELxhdqe0rjgOGhTLGVMT07zW1bnVlugkMpPBwheRAfFtEpZUMe2OCoPlzXZ91a8
KvWG53Np9qszphzBtDWsYbpnrb4xfpekcCtaCG+WFErQqsYQovNtg1OulC8megHcRoGDnpQnga71
cQckEW0MxkHNRLHYb6JGKvHhYsKlc+2y3MN1UjOeqSDWXOUJXw3R56IWTMsKVZogkSVMCU3f5AmX
c87hmXcpqqelDANOZ9rFpXcEEkgfGzIitrMOowJvbKoNP2d8RNKF9jIM7sYe5vYdMZ8bMltS32W3
HPes3u6gXud8DmmIbWDVLdkB21c5VzD9pfMLp55pVoxxDODSBy4EO1sMSpo2RhzeIoaM3z1mf58q
6um3bqazMFlAUIZA4tzCnoSmT656GTkNo2Kv9ntf57t8K4Fp0gmIC4PMPLjD2PvzCsSRAQs5VoB9
dtDeAN9xGboJe0QLZexF98hO/OwXEeoqB8JtolTlUS99SX2tixGuY+aeFhxsVOdGp8r8ozLXxdzp
08lBEZbynsokk3v3KATj4Gaebfkjl/yogaYhgwgufhIMV6WYqxFwV/RqDCWubuymoqKyB+2q/1rd
6Wp+RO4INVj9RsUN4up6Jr0Mdrb1Sr6qD5c51LrizaZoj/+8iqmCpGC8YNLIVoNvNruMPTGAj/Q9
t+P/HzKuR62A8kygbm1Hx2SPKG7XOFZm+uzWXRa8kifxWK5RgLVKT+okos/OEB/T29beOzcJ1WDn
ikkf6LeKPL33sSuBXd20u/t+3P3cn/2PY04PECTGztyff12wckdsARMdSh8VWpNKJ5Ri7DJUqowC
N4FeDidudK87d07Bi62z228hDk4ZJIYZFMP4RySlc+3wTuMIxFyg6Xd3VU9yOX07iCSiaIWNdIhK
7HxfZVxn9MQZoQHJS+Y8+aXF5nZNUc98r7RZc4hjUk7Zo2ri77l2WCgtgiUpuSsjSsjUabH3i6q8
YkvbtWeRCLRz83gN6GTc0tnD6BRFAqRsCi1c/pEIHmmzSqlVWz7S3ZsDLMwnrae+TY84uDoFsHN8
asVSL9p0Pb+VR+FDVc7zcKPf+NIFVllAkc1ckh12j4ksya9cv/jZYo4nGkyP7jHgApEqI8/j7SwK
2BHaCXQ8fHKrv++REHWB2xVpIdclYO4OOMpjpzpWr0bYKPUBhwiYXesuZQAEVRmeDbd2/COVjqei
qBYCp/uaV3obPosVyFcU4fIWFgkjBzNolXCl40gfumdCyrk5us208RPaKmIvqjZgUoBZoERpgPVf
Q8oyUNxGFgT86eE7gQO6yHAC5lV1JQlvtxqIABF4et6s/526esaYIHwPCGWAyhyQcdAk787OP7xa
nZBVOpAg6q5CvjilEyXe1omVsbw832HWYc2TEK/0x50FUyQyofmV0qZKB8hMe7WpNadz5xioJx53
oL4Ib4KMIA7nqRkQHQ1x9hYLUdK85tnIaEIjbFINwMss/QeWI7cIhN0b4NmVfzHCI1Uzqfoue9FD
TvKwpk9qdOHm6dkpoV3pV230neY1fM70eKbv9K/ni480GoKWg6AIxN6w7/G3+fg4eaLrx9v2b0Up
8tLp0K3u/JHe90gVHmeEhHmnJeG2fnSjjDmrWoz+1hiAERLmz+1oeVFjgoaxqGen/H98pZXveFe3
VPqrcxgNq90Er5DQd0EbTdpEgoQaVtumWetIW2YaXpsCogfNPINSGsqNQaL4f4ro7uoNiakYWmUQ
0t1J6biJJu4/+huCphAMHhsVqEh6idghbPcVFIb6zW1492Bk5EtOjYzOtkJSef8bDbFqm475BwF4
GjKJmnR19jkuSWaSVSAIkaOIJ9QiJGBaz6lRHL9E0TdOck9ZY045apYQjPl6gMExAG/G3A5zscRA
RAaMkkGi9P7EZoRNAmwwpHAfAsD6hSArmIdhWAzzIAXzzK9+49y7eu4BQs54PYF7WtRXIPDi4zno
kCbT75YT3xjz/I4ygR4YmqtJWN/JWFhrn8dHpGvbjynsMOfVDIoCSV5+YAqEV69hnvW/SkIpqhXa
F0GgcBr4fQaNTdHQN8vFujc6FiyOYI8G8dMbmxrrf4CAkxHPiGsbq8jEamEFm0MnSe4esJB6gNYz
Wl6hBMWLP3Pa9Tac8z+8yvyOMd+WByIIObGTjYvNPmM484olunPoM+0GgvUZYEJeYmiWZhFN6WoH
dhNaHukxvyXBy8zajtGqrtl60iPxdlWclsU/GOdwFa9k1ioO2BlCIDGLrW6XBX1XCp7l+eCFsojh
XrEgU5zr9UW4HWzA2C19yGgSQhXpFAN6agHg7xxsQU2/Vm4BRo4Iyc3m1BQVfEZdqVMoBAsX+YKE
dY51XHjO+LwQPDucSpSDqkWGJeuKzW9q1c+K9+FoLgPemst9D1g5lYoTJbCRp7srEErMZFS2wMCT
p5Y0K2HHIybfgDUqArEbl/vlDkWmjzcVnaDAl9uY6h2hChDyz7bQ3t84kyCrmMw5Yx7coS4XRiKA
quwWefDR/Wc30mX6tekawrLN2fWBJ9BHisPtoTlEB4+6gh9aKqgYmzPPDqsgfozGtTrTIRUKdvlV
pUWVNuiKQ5sbHvkeI3BnujuSH0Qmdwxx/tLsRR8sxg40rbtuiUwlCWoZMZgy9X1+2EfsdpnUQsZy
urfVzzn1W5Gv54/TmXMo/oeGs6RRBUfPxuaz85gy+BGSskxGMGS+EQZ0k84vO58O5CqccLrcRbN2
eQ+Gc5rYFi3ViV/0PneYOJwoP1KgX1WudcpruBu6NlxdqJCHtot/574KLyOhyPXs1Vg70RXcZ32x
gBwaur46Dnro+ikEq00L+WSOUZT5b5rguZtk2NcLjpmJIg5P5DlmdRKMguLrQ0OyDAd++PMR7XMR
BTvofsRX44HR/4H8TW6x8zqKZu0Xl+d/+duRZIvoTj8okI5XORbEzPauw5UajlZn80eLzWM+pkiI
4Je61+IoQ/SwHdYGrI9WAzqP/xG+nMxUWN24h1zegGnIAzrdU8afPK2TPX0m/YIL3V4ghNURWNpe
3r00PsHCbPd5ujcbY9WpVh0MUqN656Xa/rlFu4+9IZpfRBF373OdCdOouauEfYuiHle7+n4NjQvM
e1R4PGnXotZkzQXVevFwNufsaHuKFQ==
`pragma protect end_protected
