// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
QeHj3d2mVHJPyrEQ6kavjwu/nQIDwHrHP1A29IV3LN1fkMqCcKWyCl7kyIQQeeQ9d+poVY5Gh3Vx
x7KWSVEQapu4SnsHiqCAknku1YsvLMx3rbXR+RcOBSI91EPKp6w9+qzrVsPHh0SPRwLuSkGcd94j
sSFTLglZ1wsSw05PjBDW59wJpAOvrPM9hFGdJKfGix5sdPtl1LZtPohZwSjnU/w4rZ9FZxJnHur/
9doRYCvLw/lf7Y2uK06BAz/9OffpPHZbPOSf4L06xc0E8NOwkTWhbqkXUZLC6Qmd3aCtfjDw7TA9
wxEw0lXdDbF0871vscfHGnSxdTR8NWgUv1WPgg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 3056)
I8PUWwxgjWm4tI3w3vZZjgeZ4+h4ZEovSR9ahSaDSiYdOM2BuldIpxq/7hCkO4RnDkLS2GG5CSPp
6t2PogHX1efYulWDf3j6/g2PR4DNgi1EJTBS5xUqbqwLJiEGx3wORHJl7Divq2SRGYrPtTGjx8ZA
iLafVFdJoTyV3XHsCB5JOjVIHoKOn42zPwwX8txAOc812zwDWVWyqWxq2HJodW/l9R0ZfTv5Q+Jc
aTadlZkCiCfkEJigfpJL6qeg46SrMTrXJKn1yH/HDsJYUcISP65M5/AyLVg3PiXU7ZJSiReVdJG4
LPFHYCK0ox/PJc8ifdvnDOvXWUkXoSlckyULrq5FV3ycdChLLKODbpLTrMLqv0gm9874QZ0n4H8G
h/w0of8ZGUg5O6kxhWo0SztUvVSdHFYsIdCDIlO/OIW4gwHOOsxPX4UoPTXbQT/+SG0gCBF4vI1f
oe6huOcqDvMCF7Ej1ixc01bMwY9y0HFKH9GMIJGE1X4F3UODqQR1byuJ5nAvnRCdJAjcZ7jp7neI
P8fZWo1RJxCxxndggjqiTxlt/J7Zo6dKGf2kwKzu5BAMKgDjX4ZtAkho0kNfprzXI48ij3X/6gl4
taBpHWKv0t2YgEewt4Ym/VO8Tg/MgCaeD6+TNhq88dy0ejf7FiZQcp2C7/1vi8wVbSpspTze40qn
5GDsi1KELIiRZDBsrttYKLxzIC5BHZCCRPeH96g35rMujmvPLbKiHU1E5jMzIXbPdcpooxOBsBD5
QkA0VE8msYlbcfGchPZTYFTihzLvQXkH6grJTGrqzTuHAlM4SzMnlbmNOleaUrf6Ih81MP3sJ83D
wyfMyXxjhU5DIzpH8ZyZRMZieClDDtKG9SWv6HD9jxkE6rGNnBqpLp1ENHsjXbxBj0PyfZDuk9o2
E/lRvqHmNI6xSkdbSjFOUlTprhOEUD/LCLb0dFM3xMi77+5V77y0UTjzvgOzDmGcm2GJkKJzABJV
EFWcqef3FoIimkUnol+iCT765UH1+oI7YeCxr2VXiLKlVSNYCpnK8S0dFB7gwDCLdHMnnBFOcc7D
Y4qtGiP+WLMySemdcgxros+BPq9Gvbw7Sq/Gc9F9liEgEdwMOhGcLJOPws5hHLh+5rHbBQoOUUwO
LzPPk1peFmJwfCgeXlRjhzp/ET+mgL0BRcYqT/4lbIQsCSlLnwzjTiAoTXd1aMMZdFVk/RwtydJV
kqaW9I/rRFvpYhjWVUhGxT8zH0qg1d8QoMimKRLIzf9BlF766VX/AFw+J0F6cFN4ou7FQpgHL72V
9xED1VxsfJ57YZ2z3I+qtduhgwa1cJhHMSoUSvCg7H8vOlP/mG8OAH/KKUNb4Yg3oreUaQZs374Z
uIPLIYFUsdRflx228fGVdBMh3qnOOZaI4cFXT3Is9fltOWgcX3i5xzQoE9hdlhdceLNsk+uaLzz3
LPkysZJ1nNVbjxI0OUG6czpw05R+30MaPDUakRk/JQldRqww862/HR2AUCu2dcTtycAY9EvGeTBw
SyfBiIJnF1SdWjE9+01wL7B6wVUwGjkv5KnuF9JJPa84CttKR3BGpJxOfXtVZJGYAWT4H+/pOvaz
pbEME/cjl2uXnDPzz85pSNVzoAw2QRYty7zkr3q08mnGGH6OO5h0hSPpXYmG1wMU2+cvKq/U4/aE
bozvsyR+oQLdtmcZGqeQSjWkaTREm83JUxvOu7YZl0vIBy1kKr+r53qB/A7+HVGR2FT558H+thWO
JRkxZhcwB4uy/q+LXkaOVf4miQtMg6pCAEsNJt8dFoszvkKYjCpFM2fItNf/+VzOB0ZP08kihs0p
4kcNW4KWGp+38P6DAeKoiKISoObTNNJL2G1MXgYJvlDjjefnBw8GF2KXyYp1/b8DCpp9AUEJp2TU
XY1HwAbgPNxZp+0HMn247XbzDMYOkxxS79mjOTOjTBLx+DsqFpJFtGQODH+mzP7NOYltZDe7M0Ez
xthTUnQrHR5CV14+WkwAwdElvjZr+NenWseiZ/kmRoGyVwE1320LUdQMV253dAlZDJdqxr72XLy0
h0ghVpb32S5MCXB1E/a65n3PJcVAVKi4T1e8ULQrHo4FR1O35UKTacZ1eUvU2wFwITldHWzVVwQ5
agLUf0RQWzuzJzJgyFAHcKxj1AbVLGfSfy0D8FZiB6SLPxIe8+qefU3J1DsBzzPUQMn46TPZjprv
Ofd+zgaV0jGE99aEMbbb4V9RKeVV7ZzAVGOeB1uuynwM5xe+E8L5f8Ga8EJA4oQ8egn62VB8OPwc
Dmfjr7fzNN6QWnYq0ubTk+1NGZbg/xEP/vfR5cd5Pb6W6OFRORA8vtk3mUroDNkGxIDjVUkKkdL1
YkKnKQTT8jc3sR4El9axI0J+yWnecOmwlcVLemyV9Synvsb1b7szzssa4Z3ikrNaxfwhKTR+lBsk
h91gRTnEUywNFV4uP4Pqx5smORrx9/+uNLRF34eVZvOox5wygdKgzRJojLWxAanWRrvBPCfgm3SN
xqYWHFYUmQqSIAXjT1meDYfR4xsHn0SrXJxLo7cLBO43J47HXb1ShP2gkjC/nlhFmNNiPlE4hjNN
ANhCAGdKNtbEumMv6N6P+tKR6INX7D2lUKizl2b11mYTBwGcv1UI9bAoxO8ShyZeTJXfc1RlV4qs
ySTlPObNhb/RjNNFlQvKEMB+kHcjHMGgBibgzhjvB2e9EEI6UdcWsRrJslm2giYSo0TgqRZSArqa
nYB8X+dsy8+84vN/ncVusG1gWZLbO2v0302tLXuphXylTyvYik3eHfiVaQ57GJXEJ5vOK8gOTTNJ
mmOsp7X3ITFRfxSUrPsxmpUiOiHgPtgTp5/qw2jEOMfL+sWEk+4+Sm9STrgSAk9n0jYP2Pm2xaac
bXe7tboVZ+jK6SmFhCNHTNojozC2J+Y84Qc0r0t8mx5+MJZoAtytAg8Q0QCglC36n7e+oec93aIg
xeZnOPu16HtY6UDVVoyoBfFSTEv6hef44EKpuvXRBqo0f/69qZB0gAf9kr4nNLpS3JQPC2sPCd+c
XxZh56oQV2aiy2SzTeMPJVdS6C+ubv+vPq30Hl+oov3vqSjmB37NyxnMJn8T+LaoWYot0UIQPkJa
CR8Y9NdOcqCUfZk7jPJFKOH/RCBzL7T5aaROpjn31xV4Xo6R3B7YDmydK8kd/tXfT4L+YmNhdPy7
82uvtKqVJK266acewZkZdAvuJKnJYE82TxgvTar9V6GtfjPU4Aj/PdqUlsKC293MXMKduMfQZ9Ho
7KO3C3ZX92tl6yYZigZrccaFWtuIc0oCPe5IDXB4wzl9yM9yldvW0qdzGXbEEnMhPO8XdAYIvQyC
o0DXcY5ij0fzcCb+djO0CDVRdX02vsKePVboX1E0w0qYJ4lOYM7TXjaD27qnysqDeK18HYxA2lLX
yUl6kXOicbIgHixgtdWntlwBzDwSd1IqHN+JbnXAH3LxX/b4c3GTZCQWwPez9kHWzs/7kWSS7oal
p4SJq1TIFSujz704LaJZWKblaGaxMuepYebHWwi+I+YUebQm0Elpu88/6LPxCYLzju80HrKbLIBg
ZC9GTI3Rsm/LwTuCi3HEm2c00Xr+mBFZRaeafp/up64hh2JeKJV9WXv0Gcv88E08gzzjf7WLpTIK
q0VP/PwMnXLxBPqhchFOpw+z4pBc6FxkFwBpXwOjuSuSllLFe0KHe6htiuKwVwqrMFsuvVrGwb7z
sbC4EKe11z6lsK6PaM6bG7GlrsyCMn8ejHfm2CdsTKhi4o1bXni2RrGKz7vdiFftTKOvs5kxJEsQ
qrcYiWvAYnzTZAtuFLEB+M/fTCxEsURGrOwD5B5VyaRXHauFzfl6X1BQ0lV5BK6SQlhN7lQzR/cv
K70d3N8EH3+Ut4Wv8XhXSKgkGJqBE0XqHiJYbhOMEXRJIw1vmHHffqlJ2fTha+6jel+ND7ootMfR
F2ul+9V7HUe60tZvfPfWHnvMcKZQE0Z6/CEQpoDTIS7dVNjAQCuAXhvbhe87DzKZyHSU5B3yY8lF
WqleILZEIQXU5zpy6H62qeEeWZxeCn+tkV+T60JkPPNpjlw=
`pragma protect end_protected
