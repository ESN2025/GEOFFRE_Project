// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
MgwtHgeiIruV7U77mbE3vmEsIZxh1agLxk8kwoEQ0MWYY/xIK6Zt2Jpk+TmUucjKiHyV5FsJpIRZ
Y/AhAsd/cxnyu8odTyEjJDwdgklP6Gw4nCJtcHp9Gs2Pw0iJzKwU1Y2R498eEzCLexbRVp3rhx00
wjdMcqiAJ1UIgrr8Gg2aTV8E2D5qQ8gKsSmZoMJdvEYLMJux/T4JeoNyxbZI+oajCbzYJ4fgLxKx
vrcJ/LRgvKyDFfzUph0ilDiIQFf3uzoqrrlzO2m2+JYKXXAtHTDTeszJm+5/xh8TiVIsbppvGms1
rd97Jx7XdLbbuL19FTQLXwlIGnfzV5Hb3osS+g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8176)
16dzfrIOZm4YmY4ZHbHOaFI+gKUkza6QpfNfHEbd+ExvPVqcGchK/6Hts0WKfKNGqQCvUDtZdopq
pzIGpmrCal7vRtUx66V2jCY9Liw+Sqrv0myn/OHyABm7zaZfhkUlEldpfodvi/PCmtMvMKfcjpSf
Y8J09IrXv7hHpeXNBL/AUUMtRVQg76mR0R8A3bWmEijK2PsDxuOehZo/V9DXLHbFo1PMzTE11mix
yhzC9koAZWkcIYbZt0N5PQ15bPMGYQR+Jv509f4EanYmJUxtaVsYaK0pdEE1UnBmJkt92sdy37R1
Ut0mmjFWwp3cXqaB9X1NUMy2r/oA35kRu9ApG+PUKgY6EwyaRGS1jAUpVzTktSwRa7gSjpyDJXcB
sCKDh0Hl6BRMkYZc0ktA7wfI8Htr65sDcq778R85OOZTkLY+sm3QpdvTFY0CicAWewS1I2Mxbhdt
XU5sjV/AZKKe2UJq6NAYR3bgzfTLjc9FGgsILcFPLXnFgaTa6HUgif7MOkirQccHBrlcIdYbufJE
wqgCBxjhlWgwJ6Ws8dMjZbotUSyqcn6h5iiw4+clQks9bCfVWWJv3a9IGybCwdVrejRgc9GawR7y
G8uX2CDiKJcIie+S5R6Qz6e23XjfuMrCYf+8PrL9oPQZX3E2cV9tNu+pnzugpxwaKDOipJD+Y8DZ
NgK+uQELsF2EyIjLIUrZBU/PS6HomNxazWI+3F22efR5TWCHYGL1i9/ASMJfw6p8QZj5sTf6owOM
+1rnOf0yTVGKBXGNivtlb6rA8VgJzkMOCXSuMsNhB81WXHCx7ViQ4OLdt7JWRxD5MyHWd5tjf2jG
+xOzwqO152e67P8AKb20Uaw6WGjZQsmDoW+JWKH/Z4NaS09NmrTv7xJmuhVlNmRjHyDlFY5wNdPa
zMgumG8w8hCOVOdIZkSnQbrB7FMr7+MP33byq+z3DktJEwQYkJpvl32q6UWQPrjizhUS22xOQxg/
2L6Mg77Kxd0qX8Odz9bKHriEl8vy5kwsnP3aqE4I1fy7B+/1InI3IT0sdN9wHrcEA2vYwesRV3lk
4osFoBvqbEqx0nuBSLevfSrI0t7rhomwRoSLkvu+drhnaArGG2vbx3cHdWthBgKWbw6q7u+oOet7
sPRSzNU7C7E/T/9fqdRm2V885MCxzwhyG+aoSDljmBwYHDLW904zeK9YYKg8onTz7KYhNFbXaL3U
y1DB8JBJNu00aVFSoq0LGxB/6arWMnCEYI5dL6qbmsM8Nr5y/75sAn6PVSyvLDETISTwBSEdolLl
PkgMe7XYdI3GVUNPThbCeWk8SAg/9frXU9OEJfZd94/v2QotmgNS2kqePZklicTcNZ8YLI/G0vPr
SZACp9S4rYhDRzthb0GQW5uAnrdnH5uuqgGamajyIYCYXdjSgBSYHqN3c1Pn6ce+E0IpoH3i11L4
NMyD0NAb6Scih+c6q00FyHV1zxS+WloUT6UweToUc/zkCnRS+tBbcHlpOtChkiPDyc9VyhOuVkO8
Dq5uYCU7MT2mXLVfS4967nAlHCcNc5liVMOAHIdSOM/XXXNnXLF6KT6sLwCwN+XxeWmrREuCY0GA
IiC7CQnZzWCg4LGQjbpzg40eugKWpAB4fFiL7bC5ORQijhtWNqvbSl6GUf45+9YXUdEiu6bdpJXr
9d0SwXW6BOcopeuxlXtsHGtWeZwOpx67s9RPFYJzp3yz+7FCTuesZxX1m2nl+NV8Tm3lxEoW3QU8
XnnV9i+xcOKq2vzejKKHRflZ/Iicb2zts7fjzsuOxotrR/EWmWd2Vjn3WdU3bDobt8BPiSqBTyUB
1DN0hi34zTYlN8GuRUzOPZlwbvVrHh7nFZJUUfrQYQmNUDO89nm3mkmcignV3eziiBG/hKvoV8kM
FOZpzpNbqBsSZxk2BRcG78aEJPws+0bGrKh6QvbW+91X3H+daYS2Z1jUCvPdpBcSvt1L+GcZdcqq
QiPGC0uPwtEHHpJJ/Wc7PW25krq2q1FreSU8+rP/pn7UUIboE1LGiSHy4BJDV728ZZpOck/rW8/T
/lOnViY61/ou3nb4DtOtQMK8CXGjSi3xfiyzoWxeAXMYo0b/MJJEGlIj9Mvte6/zIA71jpM4C5s/
apVW+AJrCXKlWJuxhPui41v+YCo7n/wd5YXGlljGOAaypl+hnMwleb7O1MaFdpQhhK2YTu7gu6B6
vXAXDpYyoIGtaQWdIUf/6HUXrfoWjTaeGjfuhlBb9J0nIa63fjcWtR1NjKlIAfj0IzjB+/TVXz/8
Y8kfuXx1Ii9s0fbdI1kA2kK5pmpjpn97LzkfeCj9ATgWAT+CVq3YnCEoH44owbx9A9fG/eiEIbyw
wL4KlSL9yzrObGSpnxxTD6l/xImzqfR1ci+2W54dsB2U27dvUoibn95bZFgGCoZvYgFYE7oDOdAh
a/F4JN+UlQwYPiBsYFyLl2vewYa3EHhSu4vlZc0yf1Swo26GfR1GiHYknmx5AAX3PUwOcESt9LuT
rsBBaD/tONRyo1Lw+nomFSNUOWVveh0F1/9Fw39ZayY4D+wia8DTLjHF+OKQWCuE2Fga0N/81dV/
BIMCBOnkRojbW+dERlVgDLybQFcaHRi5snQh0fT/jjN5VdZ8s831F5o0h9EVz629Bno3ZiLnBQxv
IwK6B6M0l8V3HSa1nuLm/k/egkSamJfzoc0bV+5zFi3b/ClZRyBUUgg6P7E7N6CspyC/DmWshnqv
oSdJenSLOWZxODYZxLQWtmfxbTojRfBf5mm2a55rHbFgUMnpYlDIK/HNFaVeqNQ3lDRDaRJGQRXG
X2igDvv44hWcLhCMYThXMGjY4XEfpxzycjfu68zSqX7u1EYyrQfKEta59xCe7fWdaC6p1JpkYVcW
ThDeYBo9i51ULYltuZx6ThAyFFE+viNBdyWnBJX8aWkX3CyRwumkqNGT1r/HuueQdAksd3blX8eY
Qv0/IAZVkFV3nUEF5VrvWwDdxhe6RqUcwvOTzDG+kkxnPcDMtXIYuDYEOlNof97rgaVcgKi9yyAd
EmhBfwjGr3gU+QyVHvNfvCGFAz6oajAuQ9oPLhzKeaGlfKC6Fg63klFzleQy2/o58MW9K+Wg5NRO
Br25PNpwK7TgqXb5SeLw7uSDzzTzlU3dvZpNxoigT/cIMub2QFTSUaq2AXW4xzBMJXWc194afoWM
USwyxqwTOWQg0X6bFO7I5Y1ZR5CFXBSHkrTUzzyYOyP5keGit0yNZ5Sha81eyatMpNRIGvUb9FiK
Lt6N/cKH3DEEo8bVhEsidcWYLXmusHQs8EIIXW09+rB3ncUr+dlQZJhSmcNDBrNYM8hdGzdBXosS
9fWBbStg0msjOyYlY7su9PrWEiVuK0LLvDDqJGxAwahA/QhO8LnGa8F5dJ4jpIIV0DrmJf4MlGBX
XqxLHLaz9ESBd6AwOOTPsudm+Tq4Xc37jbZPzdjHc02GIZBmZeEoEnavvAHHW3Dtqg+GZeDrnEYA
XsnEfa/MqrcQLMBHVQ19EXQDpEe73m5NXXy8JnMvDYcyjWc9+s3KIzKbg2gj0bwG/ZRU3rdL5O0O
aGQu8IDKVHyzxgrQAUK3tNENHTi2tr1ssTWxiLICTI8dP3bPSrS34DlpSt0oc7rJwpH22ENP7g+v
JTqlvVZS9KFGKXgbGHSXP3KBJu++XB9GYSAPUCHc0b3yAo6KpO2Wl+f2mrXe39Mz2idIhx8Hqi+2
qVgwWfHmi5GQJY/iokbkl+qOKSBZ9NQJ2JEvIcot7oXS57uzx2NzcFOXUu1jK2ob4lJUvSa1xcDK
HT6blzY0kBp/oph81bw/XvkOKQ1lH3ncWW9uIL+InvF2i5kiNhfbdPkKJC2sfJKnAaZQdYmkqV4c
DPiJO/BIDTXwkHnhNwSzTuu4K6hjTg226Br+Tk0E+42VO68V41S4ojG8On07QcRGkXt5B5GmWbV/
R6laulprSf8dvN1iC6G322VNdFqldWKheq5Ji0+mb0Laime129SBR/DxC5lAMrK5DM5EymeZJCBo
GSY2BPIh5XzLUYgiV/Icq4wnAfdp/6/Smt0oQmry5P6V9cF5Q8C/uVxeSdO6GfmrZlwg4ru3A18m
kqngH7LeTeFi5XLRX2VpKlrI9lInQpgOT30D3xeExo0Ic8HiasU3lDP6o2JYnqhVgCK9dgV7F7rX
QCZPBa6+5nRaJqVOo+86i8YgH+u4G2DCszUWGDW17u0MSBgZtAhd4m4Jq/Z8HqC8qcoCrWjwA5Hx
wP7IKMp7wttuqUd+0R2ZWJ2UMMEqwvIMPP59FDoemAom4ErvJhx2HJ+CP6ONTQw5s62N2ZjSQwlQ
0K4gDcQT83tWY5nOHdytyLkgvMf3Hoitp6qMi1pYGxrCn2oRnyyVr4mE3GdLIByWLhtDco/OAw9K
4deiSoSk5n/Ak7Ie+MXln//v1U3upeLBtmWPYnfH96bBF0G2zuOG918zTf7ubNNa3dIZSjYKuGAH
cEgaT27zvR1NIoI3+E71hnDK7mBeRoKU0JZCQHV0YNBWh6vYnUH/TjKqm/xnKKHsbhyF903S2IJA
UrS1f+YNW56znfudAb8jSG9QbRqCuZ+biVheSW/4so9Ec9ZF15KzNCOGX6N5Nrfd6hWXefLVl0t+
KbAs1maDBgMTwWzeax3X/5iqoL5vrOG70seyqwnUYmumQ9gFr3srnvX1Nrj04GtYdATTgp1ssP28
WAd7lYl/E7p0rFAqEVA7J/3qbbYyMzuzkX9YX46k8vb+w1vmuePo3el9rH1ly2ReL4zS+uEIvv29
7BnFw790n/xfBQ6MmMw6f5mHnXVvDoca2iniIIKVKRzkrZ7Nh9vStz612dVUFr+X4PQSu8z4KTGr
BPTQS3D3JZ1/tBxj87qZPrC1oJz/41q4nEObOoIu/c3QJoFpcTE+3owvog4P3J2wl4fFN6CbusvK
jDRIxtxGm2zg+Eqc1Z2HmQTh44ZWqcfEQ9lXLBi3IyZ6TCVtMN0SZvJZ12Peh9Vtne8PpZNLF7MM
FL/v8ChoT1bLWV16eBO535lnPfGzN0F4lZvubvBWp1pyW2pmIEnfwvBR0SInJNrGxOZLjCEBlGeE
SCGoReGQIPswh7mLD7qixXu2ef5SJn1QQJB1bwel6KMReyqgGRyyHDTmRCtIiLItz8awgq8LAjld
Tzh9TT5v60BO8OlWESYU6RPSE0e4OrAc73M3DDXJ9DDhoNLV6d8qs1Ba0X6aFj6CfNXndjQubTx4
A+EUJirjNJCY1BMcqVKbIeV/37QdXEHhrHEjR26q9KniwJsqpp0Mh8yw2kSmdscvsghI4hLJFwMg
HG5SkqmP9ttuYo0wK8+B30GKRtiy0VT0ZU+NwewwIPBR466AUHznz7ECrl0l3dAB2HQLKI5Vquod
cH39zbQhAEqUiju2WMrgf9bttnaH9BrKzhevIbO8xh8uOPxiXF624QqDwXJqgclk5ul1l03TZMJp
nLO6QIlWVZT4U1bWI5bJzAMe1DfLRlCInJDdfO0AYtGBZBJSDy8t9Rrbd9+gkTG0TyOIErTkMhLj
VBmQ57LBlCyZVwIXs9yDbyEif0pxoZi5IfwnO7Gof4t9e2wouQzxF0XZqLBW7phEer4FnxWqCl3h
nyEsIuYf5/Ola75s+CI2PpsajIEevsCEtHpMr45gabRnY3h3OR5NjTBa32XIzXeHmV6+JxfyTIeY
d2NioA3mcf/1ldgbYhKHn+7w70OTtIlsrnzfKcZ2MmFMM39OxCW/BeiXgEYk8kIuK2AriGjodSaq
wcDChWxFF1vI2R1dAElAqYMDW58CAmRF/UHgsb5s1dlSVovXe09pAT4SccR7ptrja4GSUSQD0e79
U+XIifk+sM5RYYBYxOaZbf8DlTgKBul8V2wPlLXHmfJuMbRb0yKPXzWbUCA8dqRSLEe4m5Up0w4W
zMQxdrfENpux60St0AJLqR1HU8602K/qq+Zpnt38/RVWZ9gEdVy7r+Y9MpiW+yd55Ryz0Jhqdvzk
3TvGnOt4T2dW2DpYXx1GpqglyTfZUsVL/M8jXkJvfWeswanB+0NlI9GL8E0bd1KztYB2xlSNa2Wx
WXawU00Bk1CQUDuHdsn3y9HqVVGMYlX7er/4J4Ya3aYHVER/8VtQ0AVeVNycIkcSxfNOcB2tOTnL
8Asaaj+BsjQ9rhsY6DaVqcIjLeItIBsXOYZBZLY65NFnez/fgEMFFjGQAPjODuSPiN8rho8Vib9j
zZQG6/JIy9NaDbV46Vla2q5tVax4jZdbIevtMMXziSqxh7o7GaDuUFBCEc0tfaOVInZsknK/NysO
Oy67W1KjXI8uvV6LP7gWgUZl7hmRRfEsAN8lL2oG/faSFXzJjRdTKOJLIUvi19a9xXEQkNx76FDR
iXs34aN/FAtsFvoXDxM4/AjQobBvts8YI8LXdUC92u9Iu3VjfbmsXsrbFL2hi+fPlkeF0mWEndk5
hfcw0rwNASNcfXcPSAQrgrgRyqDZMD4DeXgYuUwe41EsS1ptvnjZgiA2wFUL7+o0mc2ZuwoX8Bi4
Q0LwgqDDJBFcri5fweCl01YL2XdJhqnX1rSnVSLUeKFq+aWLXyq4fsruTMC9zXt8DzW68rJycUI9
gHQ9gr7XErlP0dvhGyy1+WjnyWSVf9C1o4w8+mXil+f2bNmDxag3WagFJAupsX6DeO9IBsl36xk/
0JXofMoEZ47GfWgGiF4I99VmJ4QDWyVjux5uZ9cuMi9UIxqqfm2zS3dLKgPNWS6a67rcZeu8qUYp
CQgmadVdar05tYO/gTj8J6M8yvuF/uZHvC3ND6FNi8WI3E4ornj1VZje5mss6CphMDxVUeXaxJGd
A9fhP/DtIOVYfIE4agNUarmmki+M1qyO8zTOClzNtMgbqTE3ZKR3UJ9JCd772c5jbTMI9kK0lLeM
Pvq1ukYp/Cppq6WZHH3noubJvmscUxBj+m1jEa32N+JOQnGezODSykJeykda6XuzEEmPydU45n6F
FVawlQ9j71R6uUAEYg7KQGai5a8vcbveHnDMcVld1G0bLXkxAu9Hng/HdwWoFXdtHpQc/g6qaC9l
M8RCpdLKRnD3/jrjOrT2TDIlyQqD69JPRxSXCVGOAelEDOmNYHlTsyyU41W93uZ/vPyl4k2ydlut
sr8SydTJYw+lheGual7CAGmwuh80W9Segom1xAVOWYUlKuaoCASU7abG3IUVdrafazU6VwDxi4+9
PP9eHSr+ILOaVjaYzyOoqG+v6rchP/hR6H+0PculGZorS1LNGaaPUWadrpnqVBymdDpt/wnDiwtg
AudsiJPHHah37tZVWWqwK4HS0EKDVVaZ7uvEoVYFAQ6B5j3GOdnNXy5iNb8SkVBbDA5KCEx1TEtr
gyoUYQIAYIxl0V+jY7zaDLTdt0RDrtZOwIpclQoXS772FuYRWrq8y/YX65/nj+tEWGB+cd0qPAXF
hdLdoLc9d84bS3+ax5VHKDQliVHHjTt5CbT0q8aHYX9mtExstg4nhSK+JiOHk6G0YBOEBqgBf8r9
4VQZZ5OjFIzp5a0wwNu9354Nqe9e7tBK+QAJ15m3qbxXiv++JSTwAAwPO0D3O3CUSKlwfobyBWi4
w6Bzd94wroCn634iiJTfzBB5xYGf/TT1SofOz5PqmzkJJQdcYRGrUh5oay1jrrZxI+GgRoj7DU1m
87c8EoY9lxqCFcdqBHo80EKF1GefXyV0eHAHD3N0W81qzKHy9Gw2u6USPoegx7daJJAOWjQTm04k
E7NYjh4O4Y5S/yWKXwu6JhJY4rcbREu5sHrtUTLZrkrg0O3KKfIXl6xydZqoJGtO7je9Qu85N++q
wZ7E/KMtAYmNXcjGkhKrsTqEatjBBBXoUGYzqjJ0UdpDrtseWko8AJ4Zw7xHw3hqGwX96swwRKr/
0kLCKsqjhdlWgnaJG91a8d7abt2+pe2S7qQjLYSPZYZn1+/iAQMtJunU6NqAo2zbalukmyAPQGRp
QVyd+QSQ4kWg4DJ/Kl1/KU/1zVJ4RYsMJpJYMnuV/HG5b2V69tMLo3mGj+m3l5YaZDRhd8koEa3M
WP3fuYTnTeYhjPSlrnN/RHd9IMsa+qvyMhjqF5fQ6SHJ/HKWT7yRGp27kQh/64vh/FSPe8znwaH+
RHd+z//ZbVEZKjzGSOpDLAgZduu47+TPVhxabqDXVD6SKuBFeZcfUfK8F63o0saoGHMaFLtfziIO
YDEWESX7Q0xfJVXNhfDr8jzBj4K3IlqwY86JJb5tmu30DHW1PfKS7ocFkYVHr0PvoC7y3uzRNA41
viXDsbI+fKWXbrDrx8lr+scA1onnDPqnSKNXnA4QSYDBP1oStk5jBBAl3pp3tqDIFS5Dev+wdEwJ
3VlZ9YbD+EYzzwiTY/qwRUeqf+1ZNReX54dXZKpPirNFkVHjT32gJC17B/g59HrfVeIkp0QI8kyT
VCh+gCkOVSdw1wgdAFLo6jqgBrEEuFOLx3yBcPlxyJTNSmwRtSJQOtm6MxlcDW++NgAwlneX8HeL
kFM6ulk535hXNo0NkzSxf6ZjB/2PDnuLdOGcQTck2bANlr1Km9bAIlyvMAR6fl0PCHcsU6b7S9d2
8MJhGrZxSj3yfusNnc8GIBvHPF0Ias1fO1cl4llGmObYGlPl/wJaCOzRnZtk+D8cTf3zyo8UqJm8
LswrG2oHfQzmXU5OThHMip8lH07IJOMSufz9JTucXLFROeYJvcGIqNOrgFbjex7fxatxEK1bs49+
J033X9yZzwdaCX5Z6daZAFZjbhN/w/qkd/Ua8rhn/g4SwQVFOa3/s1f7cul1IyiVppmHYQOnSRfJ
XdWWHdw+SzHTEM3GEW22jGE32HhZ8K74KWiIjAejK7tC9CLmtEWrvTed1oKP2aseUf3sqP2RNuAl
s7hYB2fLpycPI5MNvrmsELJF8yLgYALVT8NBev92BnyZDD/qEEG1o+T5qcUt/SJU4QY3zroYcBlr
b3InKxLcAZqBVecSyb2TxBtZ7ctSfxwZFi8qlR+D/kdFKIsk9Rp29nTuvp2x7kwbxavGrxU70Ze6
in0Eo+97mFrK3mdlC1OKROVnhhcBAvV031Z0Az8FM6PZzTkKSJ/fkPrj0eHEVrsuOIvTdSSnuC6S
C9iW9myB2+CRlcDDhC6X3Dn3fTJiHenY16Sd0XzzE3vlGc5UFDAyj9MzPai4garE1zY4o7WvvDZn
bwofPyjFORF4V4oXja7xia8Hot1VZsq/45wKi8DHh0dEo0k9c1m1jJMGHsdf3J3vxVAIUn6/nX/r
Jdpoh/3J0fvrVlZBBGhVgTXlZl2jf2ZKpTNVVHdFD38C+XQqTZbxs5+aX1tYn/h5SJ8/iKHKZtDH
tafWbgF2kcEDBCknFU/l3b2Hzvpf1LOQeaIC6u36e4jNWTpVBOwQNh9pnLgjPjKnuIF8wru3hhy7
H+A1A8dN9dKX4wh+dQQG7ZBk9EX5j/zzkt9dHSeLLSXFqRUWkBt8nTAxcSlvWMZz4uqvCnlJMzHH
/ouzcn0yb2SHV/6Js/aJFNVsfaSyFyUf6PThRHTSqpDQf+HCuO0tDmQ68BWKhKwDXUw8EMTPtSNi
Tdg1ysbAF1/db748C/OMvrJ6rwG2qcT50CdWFVjEHVRaP932M6lXAceuEv7dAdep8RPYpi6mhuBg
TwWtzkWsWw+6OY811otzGb4Zpp8EL+C6rv0MUcEOHBLFWeK1O4kWbMubsVm5+VKU5rgSnOOfL6Lm
qS5dlTlcjEqCQqGePSFYt322/7AnD2PqC/jrjU1HIjgbgZiPm6mNpwQzLYdNw8TCZm2CJ8PFlx07
skHBifEDuw2zJ0WdE53MgnkxkeoWC6sncL+cXCmEu10Nd4k3aM3Fg7qjzxYcfQUAgbAYuFSoA7tP
BRZzzjyfBfpxXHUEgEtnE0TNcal48T97WMArsfg3iUCmpj1/veG3RCVPSZe8zi9V6HrQRObR2+z6
qnhJcIMzm0LjTRMnTIy6S3OwiEqQmyO5bOUFgEFodxrTQmfKj++BDakp5cbNdxrME3gKB/89dfPr
huIEMP3+Ptx5gUEwaYXlf8qRERET3N9DSXbpPQS1VAq9/w3hbe/Le6BhP+FeuLQ3DlwGHeBPoj1J
Q20yU0wrlJHuE0tccTy+NnT3QMPdDVP3Axoi1EPupL1INscUaoZOdzOp4kwaMZ86cNfR/iCimh1n
jchy1B2wh4XNHsaCji0lzmdGZgxGzI718chjLqqgDuV9X4LgX4ewuwopbOXlOVeU/N1BkmLKh//G
BjF/0yWGMfv8hWjVsL2/SxYg3HB19YS4ap8jXh00tnEFu5MM9kL0JZJT+pX98isyWF2yy0jBR37i
ngZKPBqtANCDT3hBxmdtTR59Ry0uveJRVGZQbsvfUc+nbRVgzBYXXv/EITFj6Po5A8gh6ZB3tjig
XOoNdLEta1MRDzN0eSzVCsuJczJs0YYAHivebDm/00BoH+yFJyzkziuuFkovxTpUzAUkQeOhtrr3
KCqkn858nhNAmUd3IgKJ5w+yZk/AclSj6iK7sK8kRXyv8ybXUl3r5fbr0jv2GVg35QGPaVnDWAZZ
xWkv29T1bbR8rC0Gmn278VY5MgguUA6LOuWxUU4+BUu6jV6HUjPoWkJBjuHcXhnP7mF1CqoxM4GI
S6gvPAqWEsczzinygS85HNpOmMOJe4UEmnZvKrVisnZUaejWlfmvA3o36oW2GjnVGUYoyU3jR7uN
0hnj58hlOXEafObpAdds30IVPHDu3mPszjijFHS7j66kRfc5h3CXRY/fafdqBbNwWDuqSXE0V8/8
J5RTABLOZHI+RDOrGhYSFpKm4HAQVomdCnkQVUJJUhvs5pdztH36soKe2TtSBy9CXUktdoQ3Rloh
iGem6Bzvip5AZWwlJU/N569Mf1einO90Cg==
`pragma protect end_protected
