// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
P0wqqsNZVNcoO1D3YaDQZlURMKqZbiR7ccNvIUUqLu9a2UBgqVSFuSKzaEI0aYwDW19jFrL8nn0f
zEcdM3tA8LT1JS0tQbCkSN9jJGyCVyy6SOmpxFQOm4c4Of/uquXr+rix77kT4Opn0n7uHN6ADang
18HwQN+Nz0cZ182f3uGS7LlEaJFNlcG//bLvTYccXsOioADdI4rntyeJ9vCaGAtr8AcSzxKTrvs5
re+lE/2WJM/oOqxbVATP0jRT2cf4sDPuEZRrMCojPCpubTJv19btgA6dOfxRzstwZLakkke5nkts
jnDPOegbx+iNtNCfwTSePXpQ/bvUbJS1n98e0A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 31536)
iNpHMTsBr7OVi3wgCX504L1GSqNHIeA6lkpSMaTIfHb/n9MPBO6DbL8NDtOJ+ocyDrr68uK6N7n7
AjICO1/kkLeTipggrC9LIQYqXAPriZ+oQU5K0yt+QZgCT6wI9Cpn2EQCZhfQQ7feabLJh/pmEjg+
DA/9WWGZ62gviP9NnNG9Z0wyAg+lcyqdxz3OxRIAZtjO/VR7DA8MIHYew+aYOOt0FePmDNPspRr1
VFMSsgXY6yQXWL1ZipwgWCaTu5HHJBKtLaAFQ3+jQtP8kOvViDC+NEmG8QhtQYwaR60331GEfvSV
t8+UGmGgYY0KaBXCoMK1X+3MyMvQm6AaWm9mA4I156fb4SHKeBguBpXo3vHM1qS0KoYzVnZxGc7/
Wrb7bjkZN4YkFyE3QnuRzPmdioIzBqcq1llmq+g9zmptygVpCR/i+JoftiVpCZYhnVx8IMG6+A7G
3I7vEHnnsF7o3PjBNeY33YIhvmKuYGroiCyCwOgK2K2GDa3f85NUpdRTRxOiedHCTOcuZXuG7cbT
6DXHMxIjpaYAfw6bmDzSx2J76NISxCZvVg1aXvxrpdgMoLQ4XNPc403+QKxEkoW6SazW9iqzCzQU
EvYa3pYpDQTMuetp9k37Woapi3D23QQ/QdEjGkWAEwp/wZEFslFchIUldeNQ1GSZjhEvbvL7C+5d
xc25X26ngLioKXZIqpIPgXCTvxI7mrCZqY7I0Aw28qivLWNkx8ndCe84dUGauFRqOX026jlnlfzd
VPFx6vhd2Ude/7QsZQIYl4NorXEnJwb4vOVYfB1CPIa0tHmnveV+tZYUH2P5iMgS6QcA8gNATGhH
Gt/J+t90IqJmf5lNG+4YU4h5rBjpoUK4DciEMMkU3ktkd7anQQTlSH7LYrTLiPxtKS8k1AQeWQA1
W6SSSBTOmMZ08FaM61DmJawLlu2aMw+THfD2h8geEg5wX7wqwQ82Cd0HTkisONG7SNDWgYExmLlV
mHIiZWkYDaCE8e2nyQDANi5z/Srl61CdJHsfWRU1Qg7MBDK3wAEwlyGruYuueNGdnN2LLds8kWA3
/kGCOjodsRKrCkqrr/7WKqzyG2FXOm+dzB4Vm1KtGtCSqvgc5MMZSVa69iMkPm95XNMYRB1cSxBs
l1JxTqYww/hyTwzVWTWHXcVtGGfv5qy67JpYObOulb+H5rvWZCPRTDtHwayXm0qu1TbTfMAB9TFT
anvRUKLAD/6iHTKLygvWJQBgC3uAMkPSkjgxwCpGo5o/7t4mcEMLdgAOpgCNe+ljgEa7Iah3PmtG
D9W2UkdZo/lavL5QpoHhW+meEYdmWbdv4ASQJUaqS4l6z+nv7Hwguq/tuUWbJ43XK4bSMeHYjMyc
LYzhxhGPpl0ZXd4+3M70crGE5dzZacUGoj6fLmsT87gJQs9R3FnXqj6mchPxMadzZ3zxJjFrpkZl
m2XJchpaoiqtX5KA8l4IHFJMJeV0oODTupQovT5jpcD+6NiESQCHbSZdKohIeQPv8J4kEboa384q
ZYDia8D5MIsxZ3ui71UafUaBwQoQYdDpyAxW6bfKwhEJ+Yya31ghGpPBUJBKJocPgDo+dBKGvFuG
5jthSAsQ0MgAsomEObtrAGeD7yslhXd+cFa7B5DPZZQ0nBZHApgmfrPuQxkXZN39ZiVz3BA6LXdU
b2MPRrbcXk+LQDjbIPo08GrRfvOZInTjjMbfAT1M6yQrjpI21xkJb6GNSETNGajcJKNIxhzZjQ0Y
STGvWqCRG4Qw2vDftWSBRa0k2ysp2GJnRyB8oWVzwTs6X2DMbHse/Dq/ENvWbvOsa4lonA0IAtfz
3IM2uE0wKsiryuZMHlj+6BgkEu6sjR7yH50dOachDQQi4gLH4KKMVsFICnfEJ8dF5PgH2lmlZSTI
/1wTj7udljFSebEWXvtXc//5m9Rk/Jqqo3025c6CFDiHLqmv7oAN3YNcqCxeq2h+G5BK4fJxGz6G
C0qOQf472YEdPwGMn7OC1PP0WPvYPqnoX7Qw/cRW1P/xgFbHlpXYr2kU44VIdXjwFHqFxWO0XMjY
enmyPCHjFTvCakcXAWW1zulNdZguJ04sW8xeLpsvR1LCjy2qb4LfecP3fZox3VktqoKKcpc4qTfJ
FH/lJKgNKF7NAkvB2F1qKYZbPz6VAH2tWa+iArY3B4uT+E0KdwI0qm3AzbbELvxU9sZNMptItmFf
6v8VtfRHHoWOmNeG6mtd7qS48O6OD6qa4H7vNelZ1DV5fl+I237xkORKCUvAVRpseJJGtJarGQJl
lobtkbIEz1+5t3gjcYGBmAX1VVPztWI4MEYC/7OPFFAjsA3vreVEIropjA9JKsbBF035Ycy0c8md
TVHbi9ucAtYe+7nX9elgVOJEnHvLkel0Z5sey1NxUEDSxFdLTZ3T/MILkcAHseZ9ceEkbW6hSLcl
m4ZwtJm3yyTGsyZ1+xCgjns1Gt8jXLXxmuUIYn1MMHEcbgq8N6rDMrxdKEpAepS3uaI08l2k+uik
Wl97AblG68YFOIhICpMVRQ0/Y/on8eGAEs7Yc07z/ItttMc5hpvwsUO3atLZHLDLr1XZ/Gm8eLWP
SVFykrtuNXXxAKCZf5ivYwFgxpbxZ8DFy7BTwHTusmgSwz1SUf1eVypbpe5MavmuJ8Z6VtbJ53uB
cKJZ1UDK+0Vz75mghZp9TM/JGe/pcn7WW5DibI0vhah2VIIwToauLi/oJwT+aVapMZbpu3cFoFQG
AUT0gyaKAjDWaHOGpOxYvyLSdnydWkdZ3zAMXF8K4hb1vZU40ikZTtN6MBFIQOCnQoilu1TLXQjP
0hsuA0Go1yfDT6RsFuml6+gab1oB2xMRSS9P7ELCHPVk6dsqaJcl136rkOOomJhKqO9sQN72Scg1
llmPfK/KhFtgKst+uRZly8VdIPGjl9vFaSqa5diIO5TIPpHToy70GouSzOHC6N86KToqWWezRcRX
4Eu5+dqNwbZy17Pae4Khz6TFRCGi8Fxx37S5Pe69nRIfnVdtjvI8MsgUags8b4/8enF9KguTzi8/
ZbVBqHjljHTUS96PwcSHTLtlW0gc6t+ngv++BhUzZqcKdhFIvrDYlUg3TfC2xqyWpe5O6wD2z5YU
6HinvoaZ+SBsF6q5mAYRDD+uRcmeDhXFevHrWdgRykPnmpNaSm9DkIVa6//y3hYbyM5wDBDkns0B
klHmScyvXYXFazINhkTLzwH4dsoAtP/8Lme8B9dv6YIUkESEuTYaCWIhjnOC6keDlpCwbfsdfPFK
j4jVq0b7xtJFBS+aHzGnuTVl6bwb3qs2yrtPYAE98b995gxw1KGeWvSltS9yKrYfZFtsmDSjbGhd
kt0oHESyZa/kgz2wZvfK6DYs+2amh18Tua6VTijyTTFK9u9IURehJ8Lyc4gJbLY3PDG1ijZgQudu
dRUHbfFCSI7uDm7FSJV23Q24K83YvxajdX42jISAf3k893xIE/715/dwrd/6wckedqSxPZuTeowO
jM5AIWcFq83af4585LSN+aXoQgCnvsqCWdU64AU7+/dPoh23Vxse22CA7hZ9OH/WCz9j9aa/sgQ6
Y21bJwkyVtXjE1GPnWrWxXXrXv+cieLjeAl2FdSRpNEtqmltlFmoGufp6oIdZPCHdeYAvLKsJYYA
UbMJzz5hfDHrxc2g4E7/Ssddo27rg9iIRGDXEbX3wvWBrj7jOVI8OMmJYRRE3VI2cusetaQobSuy
Jf6UYRk4FfgRZQc0dH4RmRms68TdBiMcTDF+xz+t7Z5glK6cZ5aoFlXME2/jG/rraA5lsqaZBIX+
Ljol2vA/FJ50aZsUl/o22v169So8D2J0gh4nEDMUvh3xObELlqCCOPyQT30XskBsoSUTHYsc/iBZ
Q0+Vy/dMAsPej25DfHLOvoyMrzsEBiip+0xshXhi7DdX7m4wuQM0JTd88n51PwB6TyWJDeAI6Ozh
zb2TVkvYCkEJa6ROv7TmsPtjhARCU+A8cMGiuVBOssh2pTuu9iyA1jmTo1SsZ+BIXR6/XdT9bJDv
hYzoG4mALTvDMajuCRJ4qhzt18IJkmukmWA6EyOr/bN/CFlX2EF10KysmG2tsN3TvQU73WhND9W9
77SDQQfcfXjqa+l19t+VK9geKIHISU3jtwlTjV04mmXoHkPhFzc+eyKEUhcIK1wEbi1NF/KoVJ1g
pP1k/Xpy5dzbN4bumX67Hh46NnjTsKUaTsiNZT/+rGBiBsQlfc+RVgnkcN95oCIygf5DJO9KaU25
9VrArcNDQUY0+Ente37hCG1f3MEd1aLyT7XUz6zPpghxEoohSywX7890z1AgecCr5xL8PUs8oBYV
4OXLPvYzQpoBoOmkEoEXCvgpnnPPy1ImVw54vyqBozNQWCPAB81K/IhQpxFoSg4VBhwdwcR/kU64
0Ba1mPTPNSSnun6qhkrsrYkcRv0z66mY6xBkh3DwF26CNcwjkJxQr6kU1+m+8jBT+TP576HGMBFE
TyYGMxgZ2xdSQA8sQYWL6mULz1YzixfNTAab4qi7JsLT2rkLZjKeGUKDg9uWz2iowZaXZRS81RFY
mOEaMvGtvBd4YOtfkRHfQ2+Xfh1SJ4CrW8YrPEq29HwvLX4oVuU0lY0UPBfacnyv+r+PrFpffLL/
rqfCuWOW2X+3uLv4+rLeeJiYa6rWfBBJzj9KbpbhgQ2MaMrT6X+LA2Ebw4pbfJ356Q2EDK7SJYUI
j30EdpcK47LDTaVqH++0kkM3IQFZzNFVHjUWNXamWV+Fz+1O91Md1jL42sfQXzbVHm52aw/Frz3x
fPOROeIup2hb+x4+w/EiyaAN7fWKVLZIngIlNy3yruKy3OH1T6pwX7vEh9qqtBVtZw2CArBx/xcu
L+pBY7SX5HaGUjjfbGp0NJyIk72sIdi1UgZ9UKPoPrrQkSOZ7rw4k54SAzw0/DC96Arg21mkKZJL
DA3aAvL5OsYCE1J83+Y1F5O3ntbyQXQb9DvAvqFSvHaJe1O6SqBaRkN8Fupq9cKRdkHKpg6VeO+Y
qQijV38e5CmJdcal23i5B2J++P8tkEDbZ4rV4plGAQfI/A94W6qOUMNhsiR9jcp9Zp6uovc7/uOt
600gWhWruPTz5IE4mmX01LqsP/lrkcYS9JPwLIV5qCtqQZ0EaPSV2yoo7nb25QHC8h9b9oTuEdRd
QVg7Ld6y7Ze618bZgL4BJzZAEslZpDmuFMLJNNixr5fXZvyxRJP9h26+1xvrKbcpySQxko2rF8o3
JENK+rOUHwm535ZcL+0AEBZ58bHHM9fVn3fjvnMR/8GIpsmabnt/H/pR3J2aaf0dWw48OWh82nfT
5C51XuqLmDKg8IxkdlV/dMnxcPu3tifDTGFzUE3ifo5jDo6hLn/eyLtCDT3N48ex/h6kEhtU9x2m
dOJfMwfHeQDGlssjAGp85PeUMuRchTtKm2AtjeubWr5CGXWq1CaLFmljRwnJTwThdCxrCAHU2aPB
loQfVJT+Qrthh4LNNu7d/37DT2+926DoBJsNRBuZfu1uzR1TPH+NusIfia30+RneO0My9jnLzmch
8voCXOMj4rcc3xVXzmgFtLP/uQwRWR/gNHN9nb+6dnFJS1TeyY1uyj/qghfw5/oprHtOYQ0b5Xeo
uj8sV2qfJUCyG49ZZFkclCVaeOdBsLABVMcNzm2yxbQpINqk7m5dqtIVZ5l4e5URJoaKbiQ0qHPI
SZ9XBzBnPrgMo+cMC1SnzdoOeOJubuOpC5h7nCYxkePm//ltx89464hDHUhJIS3pMEUqy9nY25xc
7QS1mXDwgVD84NYFTWJB/d6wSDahdFEqNtbVOXEGepWS7Gp0B6VuIyosTnTjq8N5aYpqg82EhyfH
C2bomQXpHPnXtT8tka39r4C1qMdieINxSu5hKmr4MTRjaD8UUL7XihK7a5n2YsFnpCvy4r0W7Is5
Yq9t0C0+FuNa693K7zDPWQIow7+TT1P3OSIBzw+Oa+z9j41u5CApJAbRZbc3xlWRcaplX0ei+DLH
6pmgFTTvjGcQqL0/XlY1u/C/aXZXgXr4g7xA7yZwcFlpunz+mT7vqx55UMMRQzUrywpPJAxpxM1w
SrR2d2lFj9/s4LHAVIEdIUjyuO+Vf+159BqIN5CUzXF2vy8VQkv+TPeMe51jOcp1U0KB4n3XveFV
Ots3esoA5iLUVyv0jpLJEpziCRE4T7gHz5RqC55Z6kcA+FV7VmynX26i3dcJENRZSvjOU1sk18wi
q0omKaDF6DYu7ZCXCAAC91DJp7HzDoV5PnlKXjWMfAOwmIQVe5VTySo8rRDs44VtCYWOoXieiEIX
Nky9WCjSe36T36q3tyi1gVNGzzRYHx/tewE7ISKFxl13HEp0MlrSLS9gSYfzEJvHlSPeYGlO6xvL
qUBci+BAq8BQcCw1MaazD5N/cSuZ64b/oV3KYbNtDqo7PNtwFLdgQeKHAcDxiLSGwEQlDLvWQg8l
1tZ2z8/xdLnvwZUqTAk8fzVDJLcecz1Xj3Sp5xsCfKtA6kJvoCS5bsRhghw+04EIdMx0Aadp9/dY
EiVksCvpGkQug76rjssbUt5IHtMHmRzHYZqkkgKWAqaxYbkqcMfMhuq15iSjKbUQsZkN/zAbkttd
XCBOOJzYWQvORXWaogXCyIF1RFAs0YxDU5/COry2wa1wie6/XYByOlpnYvTlp0jyg1jux5eQC19v
L6LpBiTv8PVi60HpCbYrgzAmGDIQj1yGVJCvx69bV7vMA7dMvWUL+CwhuMXVaMSx+wt9fS/IYtNt
LIX7VZCxKRnMxgfTnR3eRRRRlbJwOvGuF5loRHmIjVBc2QMUC2FnO5wKuFhIDa/29a4JRlvuNqw2
8bZCJ7zRpSPRA2m+LIl54fQmv9zs1rIeOEoMNC6Ynwb/dYasS31HpROJIM3JZbC8NofY2eaPnoGs
kQAkzUR/yfoJkOUneE//da88wrKZoCSJrsyOGjw9uymnJSm/a+c8XAYVWyH5AUQV09QBlsnKJPH6
s4Ab56OtOHUh1J6wGzNY4vWLriMTz9WCnPMEQMpardvmisnLVDYG1XX0rz3VnIygu7/YW9+EZ2Ee
alCqzl/GO4KIgZ1o5jR63H+UbuZumgcoLB2ltL4IqQvUP57ZJsvCDVVHBqC0s9LN5ROhlNhGdbqD
sZqSLjTCFh156Dt/htDTi+Yht7Ow9OBtn/lklgugzua9qcMqaC/1L8v8WDslAgvWOPwYvCM67J8v
M1hShI24lsF115F9X2wQKK9nlO7+iMF2SozHcnAs5PCGtIeJNvz02JmUVQSxp02eE3s2NvWgvd0J
rMt2BFZ/L3bN/vxXsJV9tBVebeGyLbro60P7De9m7JoR/wh35REpw/4zFJ3o00TFzkmLXl0dtjk2
vC2q4eVEg87yY7y86DM2pELjX00QPKbxmAE0Pj1nX2LaeQjuSpbiNwsCn7x0HglTIR1+/3S2DzGs
S//n8cOd4rrFZlGuRgaMrpbWxto/V9MG3UnoNhI4b6isQYb2dxtvi2bxlBi853GUYaQjYJx12xlu
fsA3fPLJFp+q3VUsoo/hDPSzkTe1PGlxsonIiViKGH1fMfUqfJ+F/i8wUrdqXX3QN5Rb7nISBLZt
okjMWwYKDK+a9o3JWhh7YrHMPf9B5M7Up/P0ur+R2CMVmf36sRjTgsFyFwUWI5ppJAn0vvHU6QWq
dKl+rBlJCmZC4a7mcLazTnE+ERs+Qg1lTEn41suefGQIxfcN/fqWptWyjMb3TtyO0HNlHPuZxVbK
ucQUMSaGnuQeXZtBGYLvIStE7L0vvcZRLg1qLWVmyYgXr3VIpZ41u3cm4nQHR4dbCmMjNBa5BhOZ
jwf5LWzqv8th+DMlS6ZZsA22qAmJBehSPhr+ikkF9oxYJ53jZFPB+kKW66c2wWYxGR5Y8XLVSfbR
j1HXqcqGgxQb0YDlsE7pYhQzVmdHhjMRJd77uD2jSwdrmBiUDBfRDFNiz93LINPuxG+jwKEgOe5h
vC1GtWeUrYOpn3/eNJTRo6xbmd+ohbKPgQU/2IqJvMkEehT5WYswvjw7fDLmR37LJtxla1dHdtVH
qSL7Yq3xVLnKeKy2QI7iY8xBJOmSv77l46Z9trkI3KNW+9UKvhnIrcuIcxBnSbp5DHrO5GYoBahN
iuRfutGAxSCNoK4WwG6dG5xP2FM46wl4H4GKfL7B+C9all2V6Gu426AqvQAX33AN+FervN8iZcKD
kNwRvxx2gL1GaeeimkEMVz7HNkgEusrOh9C8+9VjrVE4btny2B9YZ/xPV+SBVDHC6GNQMHg11zeS
mdkHThI1sb67RRlN2rZNpZrKxzb4h4XD8WRqqDA1HZyU00GaEGFYHYv+RqrY9gE9XFDHGHOYx03z
Kk7SAzKmmQJHdVsJ30EEZEw1kvolVcKlbWUNI1Us10UieZeps2CUhQw7AlMhpd24jR+2ocQzadV0
seDBWWpBI/QpjPHSTQmoczix4qxofrxxPi6rKAxJPUzErTFcWnUxYW/VT3R7T1XXQOS1KevrpoHE
WL3ab0qXmsJXimFrryVgnw/4P4qLECtONFhWPklj/4MofPtjSYpx56b6/Br9LpYd6l7cg99bukjR
4nNngpy/MJzpvDZ5wo/aU6q/59ZbBy+GSclAB7W1qi3y7iYA8S5nN/XGXlklfSULq+JAL4urcuux
mlN+oWJbQzWRG1+Yn50mpBuE8xzlXt+xsmL8uZ3YElvwY+jiFMewJYUzIDTAXqbMwnTJMjQgHZOx
hhc4ztkuIwAx58oA2Ihy5XO/pZA7VgMKANcaiqNoHl+oS3zcj6kZI+HxYCXBqMFPwROOMVpnU1QK
mCCiywl7sfiQlCvwFxswK8Md/x2lEgVkAQO8iZyxGWo9bOAIEMLJQR8VMBOVGjnW+sMW/q2JPZwk
IxGzcfbW5FxgHZgaoDH3NR8jedOTi8N+5lU59c5nqEQv62WyJvHtj1oMYvHcrW372NSxqZM3mcra
svvJ14Tn/fXVyewno0+qUpfguR+Dzh9HGEYNj68D1Xehho61na0DsdGmywBVvUIw/g9JceYpSfSR
bCBL680yIKvANsEx1rZ/uas29iBsI5JvkVQMVv1IChfqXvqGkooO696Ly13mTI299YOIOIH4/21w
psHKRpBPyJwEZExXvlthrEKMu8/es9h5pRY3DqGHKqbnlT0OIUgT0bRjbSjIwQqukPdkJyZQcijn
fYpOOYcemVBcEKE1+5gWkam3dnT9UAVK7u/BAb2Hn+A/VpxKdL2GkEpd5U/viXNDEtc+gd+MSvh2
y8tkunwvpplbQayIYwV0OMWseFmWgee61lYnud33g2hU00Rmsfq1vCBh0FJE2+JbmnzrFZJQVf0b
es5jRs4YOXy4mF7jfLVSii5dgRdKCd9MFcOv+yVfJONNCwvD4yIOmuzr9/e4EmrkeZ6/NpBEZppR
FeARA3P+03xwTGSseYFsjCLdziM48tXPPti7kI5Us+pzMNoV29bXAfOJ5kh1vaH69nlEJLozW+Mh
qOkM+9zqKjZukH1isZ5ax1bW8iHegetOcMVW0EiXHXzQ3aQ/2zdi0FvcN4bFKNgk0J274KvY0zD3
RefCXDKgyRA4c5Ix14OaJw2n5yz9f1/J4Ac2PRJBeQcf93aS17r0KjTAiC3tkXegqGB077tAbXax
Qc5QN9ulrg967tJaPSA6ZwRLBJF76o5uuij8KEAI66x/b9tMCmCbUg/DFPmiP9siOnhwX8YJJA9P
E7FPsaDgbMvjDjKtP8uj5wkeMHOqqmpoGCBotkqXGYkNmJQndZlQYOKyBzQeYwvw7jQtKhC8QLTH
E9Z//m0n+4wu3OYmx+5Bq+Z5eSsO6lIJrP0AVtmbIYTCNdcc4aE2GRtfJqDIWKgTQ2UhCeyZy+Cy
QCl0ji80rVIfDmcLuhWArPd4QomNPfA3eAWYVpG2NJZVf0r5oKmdTWd4ymnVzxPfNMG+BjJoyFxg
SNDOBkbJg3wFGdcnv0DhD451mNSYrGVj2WrEcoobBoItrrH1ThbWU+i11oygOLMYEy5RT+X7N1vO
l5gLo1XLy2nfpN82osnXIZjubpkBJ8UxmY1tS4u3pLiNFfT0vXkz0GvYOjTJrYyD0llomLnoFhs/
ijk0EFTs3X5S88Cas+ov7ZI0SZJw83DjhND1YGW0eSn9NiXtGUlHvrOYceiT7kNysHA4JyV5Gsx9
VUa20SwBFEuO/noAG6ks1fUgv+H+qBIdTfaOHRJXypmdLU8+CbkOj2KaTM+etsDCw1kqSVZIIfus
pQ0JnqFdae3U92ZkrwkgdbxcIuAGB796gMiXfXl7TY5KXaT/ec0YOyBJuv0kovcM+OZp7VvdbIWA
RaNpvsUgB1AqmcPhZizpS90g8Ttp0J9xjJrtQ00reR492hzV2yWyC4YTPXpkcJTn0iHaNL8+Ck8+
bZJ2TrOQxWLF34ijkaJhXXopG6JzfrtIFC7GTrrMokZ65n15y05e5iDhxnyS3WXwETdaOzFF3jGd
vaYyt7YI3SDCnIkS+lIUQPHvoff5qdQfZSt4yvhX6LW8+IhVTy4R2juD0GLZkp8bDbpRihZySt4m
bMHCmJGGkSSdjYc2V/nWOWB4VppzI0xZCyX8KRaqB44PBs8ppld5vSFu6a7QwYpdg01qw6Vq6y6i
0vBNmlAdEJCochX4vhTYLh9eLK/4zOOHwvWhmq3l/yXxF7PQjUCE2phSdP+yigDk2z+7j05WDzwQ
XMtFcSWEvRfOOjPx53v1tF+uR2uq02sfwgv7Q6Cn7WyD/D3S2rC2uV9wYqeEFJ6OibD47pJASn/r
7jRrnaAZyWl/nA1N75B/reetHIE08LI5MO6pOKEO3eRFpdcKo4w5N46B0U5cOFvSnu/tA3r9ZFk/
Omzffq4Jx8LqyjH/Dke8sb53NkBU8pB+srY7w+rRQwZvrbkFtDTH9Ze9v8OR48aI4sbNcMlSKNAh
L5Nv40SuDvvQJt7qxqQNc8ui2BhSuTMdjmaE0O0Q86OT68S1ycKJeyF89AGUaXckmDZGldJaRRBP
7oFflZ4zY5Sm7Jax45fktyh7ICYH6gz5+GJUIxEg6r1dHbB6tmtPH7JvhHZK7VPbcvVzJrAa8gW/
vbkjeIv2DsvJCv5yc4CZm60jv16z7RmNMY+6A/q/WiskJ+6lFT66i/rm+oSab+zdge99fTQW07sh
n1S4laxtZXYcT1ljR77KB0nD5upFt0dX5sHHbZED61m2Cel6XniRNcHpa5muKco2FP8OxKgEFwbc
ry2jequ2qERukOjqcAuHSGsfEZ3rnNBt7+nOXWzH1jvZ5qxze8rID58V7uNz2+v+LtiHvUmKjw5N
H9JwrwaG3Qur1asNRJS8aG1nLG4pvrMCr8GlFytcN/ZHpIsU2H0AcIWtH80YqcU0cBjniGU533oW
1iB08JcdVWFJxs9Y0TEtbDiUKUdE0sM1NJADHUK6e//MURTW1ylljBtb8qt8sDq+mfnjH5wIbTm9
dNQ1nRIFlaiwXR8rMoFgOswSmZwDYF57A/Naio1wmJAJFLh9IfdIotkLAAgBNPUIuDMMnGCW3BVg
cJ8x4V+uF4MDrL0nhgJuT3BTh/ifaEuL2Nhd5PuaM89dYfCL+uHuF0cCjKdVw+ICe3bZorKs7Yxr
VIcHFGVjq7CqRyxsgzhKHjwDV8mkoJ628PWNzqYItLAaaxPIYrRG8EPF6HcQr72JUgkd0YCPUhZa
9FKaVvdkjLeQQsNYZ7KVuMyJ8BJIML19LF4dpfwREY284GbrFSQoJ45KfEd4f4kRmHQZeiQqYoCm
0P+yB0qceVeiP7VeLQzeUQcEBdzOS8UmBsDTHbTzj8IjNpGZGtTol41rdxwT4afdI7rjug4BZEZl
XAUKg+foOi4egkr6kCRKCFitwu4SPPlEcl0cyj2RsrhBF9cQW56hahmDqmNdTe72h7koTHw6psV0
7Pe7eYAbn6Q5eXdHi5BWbpGV7pJJe1RTESkucbFLEH3IRug5Q27zZbTOn1mFk9IjkNuXolRT7+Du
wep1Uz9W4B9Xm7RRr3bO91E8GY6QNFxKGQlss7MGD2i0wMWBrAh61YuQgI0du8yAmfZnpcCmsnUA
kVjvoCPiTIvwJE5T6siwD7oa/LauUBaeGFrdDDOSHatprjksLux5Hngi65VrFkLY0yry8in0Cxnh
nL0Ck7GuDpQ02cXBZyykxzTGMENhBK5WVCJIXjvzdBDgTxIwcwElICC0Wj4OHPtC8sCy5wa9nBOd
0H3y0wQLKXLUo9MDyT1uciB7nqjISjjC45oTpmaw4YTuaGQ9MUTVKrYxfkkIc+8/4DPp6mTGaBuT
tfZYRSxSiBXJF8JEj3ooJF/l3q5y9xLcr0b2eZq7JZ0cqR6seIdO1Q41vzIMcGB/Jebj34jJSN36
SR+xSbIsjocn7iCFO38cFuxOj/X9ewyIeKZ54xMC8lC2N12/8oNuVJKqY1q8hGS+OwVSbqfkS2zY
b+zCU5n4jBqdrNYfj3/N9JnF2IZjuo8SYSL5h2CMaaJwYRjFAl0HpNPBUmYx1i0Mvb4aqGm0Bss2
a+f7q1n/ChfGK8IOIdkyjh/5s5LMHRFONrvNXvIr3BOsVQTsKflsMPRpfeULxBx8l9O3EDruNMQg
yuqJHXvhVjB9XxcwoVzyNtZqyRMe8tGiTCXtnDJjY/F7j2iEnkzqQLA+Tl7dcoq67rzzKMzW96pC
S88KC+6vvYVexBV2Jdzj47gTeY4EwqxK4R1xcr7YsvUt7i3ct0v7WfVXduXh/EjKkegDw+VCT4jh
EEfW4ZWKEeHouH89+NMHz1+nhPthBxjT95N37h97F4SIbGlk4da5+WjbGCbLPfoDmSIUgcgI9USF
ZGQJNmmWNk71Po1w8QuMGEDN43scj14s1jXnfvLSZpyV4DZj1yT88GhbhHJXHrVhmM45hMOn+1B0
c+Wtd8utZtGW1pChHpLzEU0xLv7qLLM1h4motfQSe+jNfC75ptKYMzwZ0jnqIlVYwhbZK/AIU/9y
0n3vBH8s16XynJTqUbNq9/a1n+3eCxe+eO6aS263nqtMbAMX83ERup+tl0t6vHlQgydVLpgbNqkQ
V/f52/tQB8qnHg8F0p5F5+OnGOP7bpWE9TGgxZqIhreIxEXxjkwW7fn+UI9xIlPhgx/O0rFf1RmJ
nkel20cdeuSm5tH9nOiPQQSMbvP1you9wL1jb8XAItjIVzwCbSCDCri9M+bkNuPMKqiN+OO0YG8V
3Ns4tldLo/mhYbFDvAp8ANBQYDeMnndskeSzdUa8HX3pfV0yku4kCJV9A+CR2UPzXMY3Chh2zjVy
9ZasSHxVLdmihTJT8TAFS46OsW74OFoOW5alD3LhlB8HyKJXBy4ZkvtXSEB5PAkrfWX1S1MDApAb
yiCOVcAjhQktJQZmUV3xjs14xdDugkvRuLxs/zFOJ90tEMHkhVIqGFhPLaZ1wAK6ei7H+gIW8H++
U1hKUPoSdV7vLE7iDONd4oATZM/6JydTwPEbPVmi8us6ApTd96xrKlq2hpulue7XOZ24qJsepw0n
y1zFBy1xMmX+dzIT/n/j8fC0rk+jO/CpJ2qvHpA5afJ2vXLu8pc4VmFB4j1LGJVXUlsQeuUlGMGb
6vrJM4sZA9b4lvhNBoWFq9cGP5XlUC/0PDyzKV6jd6M0BD6RQGd3s18paxYkTx7JfAuWtOgz3ffA
mHAMq+/BFsc+IsgLMVkIIJQNY6xzyiyc8M8LtTUpArCrJhDA3HUZw9nHg2LyddFcZZlXXHC0eB1h
uFhATv/4ZPUKmEGvLHryUgo7ZJ2dnbCLEvtl9LdDMoHJFliCGwU3wv8ovW5bjatBYgqcPNAztBg+
5ltEIMwfHSYZFx4qsemis4aG5dYaIRuC7n8MjW8J28GpzwuxUwk9GiimXBrUcNW5zHdf4xPNl6wB
9S/xnGvgJCYMkEkxokbpQqFcQIesA7r3zfT3KZEtF6GoOk0JL5tGIbnng+dUfjQvFarXOOs6LatL
CyGXAF+H7XqM/gG/gtdsQm/lAvfx7mZrgZUn8zoGcfE332MU5Qz7PYWTOYqgWfK2OE6AwAP8gfjy
nGsAszHnFy6hHUhTUel1HumvOQ8TXiealHIf9izgzvRPxMlOcJcs8qcgoc2mtwBK3UaA/lcn7boB
8244X0TlEBnecH2pKNyd/Jbg0QEfxa6GXN2f879lvFzzUENGLcH7nisyhHcyDJjnW60IZ1icHe8m
eyHotmEvN0UVCb/eSg+WRKSk3Vb+Vg607CQyQzj1icOc9bTqC3bDSjO5Z+kWObVUBVAfQIhcCq5W
RBWs4r6fXJijOo3eNKG1xG65l3giFglOvVTnEDRWTjkiv/5Zh6jSSSDmUOoynU8XUnTy55KA/TvZ
GIMQCf98a2GVQ1F9+JM2awhFUhX9a8R0Jk95gGMTAUYU8lFCyywOxD5VtnJ2pklnD/RPSF4Mo4+b
HkySXnK6FhH3WdpMPEXfyvT3OkIPZp4+3H8sA0SzpnjNVMQNw9SE7Aa0YC9q12FyHHnQPKUZzMn4
0OecvlNw7OHA9x81NowoUOeDs9/hCmKAAH8Q1uxi+lP8neUF6smWfUalzWg6XNt5ipMg8fn1/JNW
KcmgfDGSA5DX/zfcynHQ4JiSmL2NFDHHPVjATph9Tpd7msB+MRpsymgoqWEjRggESQoIT55KwTnJ
XNOM9rrKrjr6o9sDo4B7bFpo/dqLPRDZqx0xTgTGjkJnk14M6t7PiVBCtn3pIlK8VNBIy+uwVC1H
OPdcx/3Tjm8OYxdulrOgBOsj/AaRdT/vXa2oEi8zns2lMn18dEJ808q5NFa/hf+n2VqEcEMh9HRu
gpbAtkhzWENf5cXSIt4XLLNcL5mBnT2GOM1AUSxMX7H4ppEr4LGCRs60X0ZOviQyXvNDhAKrDyAD
deXsQ99ln3iOeDCTYiV7LU77DItnKO6I2BjxmeixkHqSxmK9liFnZj2aL4J+R5e/iNFqWt+riJIC
lY/zGkdgpb0OzXifYJx+TUIriR+rs1VXllMlOwrK7qF8SMdgrOXwpOAAJgn7tk+EYiC5cmBDoIhz
0/AA4wGMrPOsEeITiiWKAG51K4QH5wLwSzypDBitdxwTuw01KS7ZcyyZt0hMwb5Mpq3FeviM9O/G
A9+fCFLKn0Rb38s+YRdO5QT3judOiRevnY/rIjXJi0PTCJG0W6ewWD9ghJERC73r4mYQrQ0924hN
hAZrkwvMntD46nJq3bQs7EqXnBvxrVRGBXwAVYyiGl0ucThxnHGYYW79ti0/HRZxBkVThn9+gArl
st3xsIuMLr5Kuph6lJLi7LMbTT3EAo3NxOb9BtEKM705BxCjHi997ETydpkecCPtbu6WRqM7XZ9v
xmuCN0e3jAP0cge0ikasrN6lGOENmDCKLHz28WFPRrc2n5MQUi+0h+epiFtxeBUPURBiyfHJc+28
HEuaEBNAIwPgwn244RbpzIzJr1p/tWuaky8p6b/8C67LctYgFNFv9CytrOrqgAGL/FwJUd4fLHZf
1MV8eTaUAuc7zPfYxwkeI3dNzA3tabtHu3B3MHg1FFUimL61qVGX/4SE7QXMHEhrFpUSKG3X9lAo
XNIUdCDdNnb/MrHxVl2bbCzPkDKYn+6DhM7vAVS89xqWk7gOJjMQ72Rj/S2lveW1Yb2MbXedSHNd
wtFOTFztbsEZfbU2YsugrOn0xXz8leZmrJXglbgTe/ASZv6wo9UsY4VR26jCFOOAIyYVDX6/e6ma
MkRd0PKsdrxs7Q5IwQ/TSplo5TGgAVhG4cYuYaIitOan2OhkJ8fbFuyYxm5Ad1vJtIB8CSw8t6qh
IrzQCP3cCgDv2pOpBK++rfcgN5B5wLMz74UDj8uqGzAl0HuSNEF9BZxAvpFfW3nqUCMuIeFMplaP
4WY9jfjIgEaL9TcxZgtTJ/ssSt7CnFyWFEEVrya+hCNimJj4XmddY53NE0xldHv1hRhwqfK8KULo
E35DX6lflz4lwhc+ArDlQLO45nF0TFX3+R6lusS5TaUwgo6vIRnhUmv6HWoFfE/s9wN5tARyHwPf
9fkvNZeANf3Qi54jQDGZNUuT0JI78xtqcpWTn8l3hE2Oqk78q7iz8akND5OgROxdeXOeOjvlLhbt
0ZAZTi5DMvbkiinkn6yMeERnjK0onNuy7wCBkwTCrH7S5I9Ch93ZvrStSlaCnOFHnceSeYBfAEmU
BrLof/zqR7OtsuHP+TqaY9CtxhjqYRnqxvRUUW0+763oirA0CYjZjt7vWDykE//WXYW+XfIW34TS
/mvZ1yEA8DzvtoaT2LE8lRbiwY/75Zm1q59o1sj3TWayXYGk9Ne58cZ24MvklKF85QTj8aEup09c
1ERgSm40XJC29hXFurChHI2y9qwifybaAfN4FsKm56SbNU8+Ck8knkzseiDkfREy84STf4+Ss27w
NPiabEOhPiaFOmsGbDJJn5OB0qVL8ailZ37lpw2w2P7qkyTfjWd1v0p0CG7dkbgdNRh97GX5FqE3
hUMxrCIeSKnzl9sOOXIrBvXlGHNap8OYOWFzlGMJFTHwBlT7DxnPWKijw934Jhh9XXgwOAiAgRRs
l+xAMDBwc8Wjwsj7dDqUuYtTR/q3f/DIaY0D+jwX7ticWKd1dmaSLtnkx1biEctdo28VMyg9ydjM
vTOhx2vjmJfn0xrbTSjo7rMdhhsk2RWaE3x7DLt/R5R99buFZ7v0FGSyUN1RtY23K9r5uf2Q9hm7
oy0x5I0ghq/IVmbQ5HzjhhO86Q5Veeoygm1HBNk5k+kod0oEElMC87Ops8atng5UO/LQruliOgkS
KNvSS00eOPMb84TvV8RcOBneKKQADAMVIPFCxAAMN9D5Xcd6eKE9r+1HI0Ng13PtS2gj3UnHexvX
yQS4axVtGErTXkPw2H6YQfj3U72r+CjnyQblHM4K+afYw3KaaZhAPk1RUjQKazrBieEFC1B2ZXop
Ugd+LP6o2Ota6gbhGJyRmsP+F5z0Dh8Th7v8soBzT2A+folaWyAN47vr8j+U+1HXkYc2fzgSO6Cf
igkHsbrY62xkoVHvy2FEEAG9he/wUct83rLsCgXWj9SzC5QgnuHyJbJq4jGpq4qj3Y1mV2DmKMzs
A/S0rxK0xZP6lGFABziqQ2/w65iaNLL1sCKKtPiKdVxhkC/Kjo7EKk6wWMbF8HXHYKiKTIlrFroN
JHgZCH21H7RtPK6W1pnvO5LjRVF6gVkIJwK0SzgSMfghPCNqsmEt2VdCx21MhEp3Z8WEgbZmF84V
tMo/SBTRKlbmVdnu56KfCl6HNuq8H240UqPgUhXTfUYHzotVv2oeO2GejU37r5clequ+nIYmbabY
h/mTAceHZgiiGM2296psfu26wTpj5PCwpn9ohL8cYeFjlxYQHfQUlIQNh1gdM1lrXyoQvfx/+e/e
xZVC2w4mVLuJDj6mTtkD+8pfiPnAyQieRrH9Q95gfG3Y72cBQghh4u24lY1hzHqdvRQ2dEPhSXxq
wGUaRUxz7JiVtqtUw3crj3fAH1cCggfcG8hLnT7xMdmgr88R3CCNUSIaAGlJA6nSuGWsNEQ9B1JU
4f80mfzCfbg9Bl2vqVLF3X9ki9cmDze13Tcy3H/1f+mFxMdq1EoEArr2WJTsADuIirYKvJUcd1sy
hFhqEZlyRQp/lfH8w3x+8VGJGji8ksNIxzInraVYPB/4Dba6Ftq0kaX1ygBlMO1Wfu+T4S9YBquh
G+X3qOJ0xbnp7x8mR+1yODLPJqR5l6TDtc0Km0+gbmdEDdWxTMvRHjrvW+1wA8d6xSeB6SgMjgoi
+r2Cxz5BgKmStxoyJDOrfC62zTCFLuC8WuUxnClD9qYg8ZgjqOhlXT3KdwCaZni2fawrbUzGuki6
AXD4ReGpgvyMAQHBrtaVSecxZuJSnXm0N/7PZSuU6dfz/ImJ5eicSGLD0S1EmbjImYWIH9RbJ6Wd
FjBFpWO90BE1rn8WxHgm+vt5b0NIHwewYqVC25TbkzHg2BTc5bRM2mpNVO6de/uRG2pY7aOJiuJe
iG9EUx7OCtpEoa2sophLMFanmREoJotLevaq4JQJsYvMYq7NVvhRg3VpiqbKiHL0DwV8hrcdTuZe
pzfZOVsYfi8aKnRJ5kNC1x/hYmZs5iI6rieW+BwLoOqUDms1+xE9uhluYXCabXQYAHSRsezazivT
lsunK9JN2iCFhZ5BfiKh3KP7R2LZQN0j+cewt+KnOS4hNMWO3plRjo8hPD/hHG4YxV8cBuriwwzX
GbB59zckzgfTli4Wb0YugQc3ThCu3JEfimjSf0YyilvTVctPkdp9QDFJQKHtWhduboaxi+eJfrXa
GT1NrB39ugkaxiWyXZUsUsPrFaQQkQsfhfpC/wguR5ueB6xIaw7SzuL7VJhskhG2Sb2kaAZnfUD8
pVb2uV/M+bRemlDlp8FQGRQMo9yhsYv5CzbIK5Vy7V4wRsIpAXEVKX3BP2ZNF6WxGvnOIBq2jztS
uB/kixEauOzYPlGQ6BaF1m0pWOWVGCr/H08/n29PCGJExqnjMarVw/4gxFSY84lFkPBhRnsm7RRQ
r5mxGwsybxN9uMxB2y6vXIM22s1vzFXRKrJbr43iBmj0O7Wp5fahXPML3vo1nTnzdvpf9FVrqrZR
4KTqo3Kqbg7t/DrGbRWZDJkVd3xOqwyqSllHMD6Nt32If/6boJA6nAQGLdXFrmKwg+TNFapAqhQG
2O6jvgg/yGcG+u+Wv6Hu71TeiaRJ3qdujnMGmw8LoXIowvCd1v9T7ubOdq0PW+ufGbMTQrhMW0T4
leqE+xbioyHLybMG1TQAWUz80N8PAjAYnVkTpqybxz7nrYZW9fEyL2tI3ZPmTVBNN3tE16bZg/xH
zM0jaecTijmlCCDDKgqN+mjKNzPiOWsv8qOiO13fMgX4Z8yIov/vpnGgowVtw1T6GyGKsUqCE9Nk
/TpasbSb9Jm/S2DPUc+6twQxu/kv9V+KSqCCZRkQRLOcps+yGYx4hc8y8lgLCHXd01gMtP3QIxOC
IENEX0fNuJdAz8RHVDk5c/gjuikCtiXVdLV6mU9nV8XlCEoX+tJIQ+cTP6HfzsupQb6mHU99oWux
W813FyhX905AGeLPJCGt359XItwHA2difZQ7JsiLNfzCY/6xBaiwjJIsIcubSOk0nFhbY2YSmnpj
PIwU0+xu6ftRovCindnuilTV9DjL3C7JDJx18ZOZ8d8HDhpDs19Uk6p6Yd3sMlU6cVmdiQcD1wXa
SUm+TTlfGkQHRBlj3HXIpqwta0Csj+f/uxUjF/4FBwiwClHXPCaMBq3fHRsXzn1aiDZ7U76CaQR2
UI7v6LAY95/LfuuUC0bFI3gGbFKe5qkdkmL6ubgRNOUrBqnqqmUv0rj/C/0HvNY7oFeRSTWBi+9x
uUDnfA2OMTZ7UrasYloNc7w8RrS5OnecIacHkCU/SOxxn5hf44UyR65o1vjtee6KixjnbW7ZxF46
AGTRt/R82BGgyC/ccCrZ4+VoQ+qSd9BPJem080Zj1qcKLMCkakZyeUMDL1WUfxPJ7E9RLK0ouaSl
lyntP5y1MdbLkRHmmicmxmvRABf9k/IuaD6zjtQW/h9dNh1URScbstdjXwkmjchpJ9ULoM861kB3
dFO/NTL1n1k37SVDpD1XNkXZ+gnx0M59YbCWckyOyBVeW7Ho4jBwpg2Qx9nJC4suwvGaJgLPbhrD
aQDDS7ABx+lmK+NSrjEN1QFslT2oFcfi5+v1zI9Z0XsU5R1TlNk9/WEOsicycxXw4nw5CLhjKh42
no6PtZuapBL4IZNAhlXYO6PmPiB017K51OB7Ai/pntwzIvqtr6u4LxK6e0i+ab5qi2PR07sHHjK7
zBXKElaU4X2mVddiwlDAFqBUfU6zorO9SI5tCNOFiq0VnvqDJEHRUxsmG5lxfnBEGm1/RQrOlI4W
WXWFrQQ5cEE/tFErBVt7R2l10QRCyGR3vEiY61aHSoJf2r5auu1XgSFKgt1kICuhV3QZkR7hUXBs
CHkmeXXx8STuYcNpOchSqbHViPYbrHS6JvUYFqCpHbUfOFT6utmFJZx6E15xyt2drmawz4gb+T0/
1qIRB9ImNPWeL/eGcqL3dT/5Cd+JzDdVNi75sPMqyKE7nGDy4Hz5cqaGkPiPFnSPdG+sAOCyo/XD
1fXTQCf+Ol82BpX3FnY67+WME6VCR5KSBW/Glo45dUoysYKA9n0aoVwu0kH0132uLgc9dKAD5p6X
+F0Br9cOGeEiEkGVyXuqfm9G8C1VGPP6o67/BLa2q8J6y3U3aSYhPZ4yd+W0Lwa09qLvXdXfgkwT
M7n9QilDdfA7foVGu8k28wr4CFzHb0zGZYVnWClFz6UfIvSK98Keb+yj/60BmS11k2l2Jqs6J/z7
/nhPgSO23PwRdBOAd47ZSNNwJ21N994XQ4YfWXZYKQF0eLHBoZ8Cv8JbML79WPNQFgV9fN5eB2GY
sWWh5Rfx9ZiA9HV1fLhMJQh/3TDe9x0FmR02VkaxqzNlP+n0wevc3zDnnI+cgqfk3uhiRTnB8Vj4
st4YZL5Qak9RBGEi4T9jqvWS7HKSAeKyruO2QFxhvCD2NkW6dBCUWqhBBts93lgs6zOcJe8j92nX
Bz5Cn6TWDS5lHBGf7LuzhiqJqYv4+7l2FrkDRI64JUT2UCqwL8olNaBz5rfFN6EVVg/PbwCcv48u
yLxu9ptANuLf7LDCUv1QjGuKPZB2Bt3V0O5rDtJv21xoiF9mNTKQzNscDHvuD+9+ZuORSXBhjprT
+C40fQrt4DM7MmpDpiUieNgaHBSxkB8UnkLL4BxcNhtDaRCp5ocYeghAThB5CyKRI3pNvAtdzEOH
30+mYdyccRcIIzn5JK6dTEZC6jMbWIqpFjORdc0Vss+TSjOkyJkhYSni1SuECuqH8n/CBztkakBG
eKauaAL54RHfBJSXjLCOOwD7PVWsKZ07iZLbwTPppfJaGvFT65kJwRRNwypvVTEQPEfvgiPsBvEq
wFwklZG3UMa/wtHgSY2BdXhjhEvnuXdjnEwhJqP9vGzg9MKBJRpXwdnFxHL6wVcH+GgQgKUzqZCL
maDClpXGLADS/ndDaB7+c/34aBU294m7rvrKggYd0lEFHsWVaULN+js3UQO8S4FCy6pa3W4C14WF
4vxpoe5c6AB+Elf85prcfwee62rJOg9V3BIMhB+L7h50GpTmYxCTx75P3T9ZCoW5gWcRvg4wBChm
n305K27/5PodL/z0835snrcd4FlHwwEcu+B0v/gPhAcBjFu81PLX6CSEkUukN5x+XMs/bmJ7Guic
0eDIzAVapYUdUeqaSV0V+OV9pBFEt6/9VKaR1MX8ZwwxSqQVNw5J4y36gsKJqWtq2wvA/dYLY9oj
2FvM/j0rrokLrzss5iCLcypt9KBzDwqpgNGmI9LTjnUptiWIw4FAd8Q/gd9VtrOdwc29r7tXaxw0
aI733KzYGKSKVcOStqWzekkdbDOC3Q/6oBYZdPp57FoUsuUgLp1Ofz9iVcYc/IoIpZa0gvG+sZX1
tdZgiDfaqbSZyAGSCIXsBitawh7AjOtx35/9VPCXDAV58LJuPOw2mcqBxCZF+tT0vP1X7q7NWuxx
uV5oUdx2eSuozH1GDj33GDF1nAHGd0WeG7msgo0PynkLeNRGlEKZRwXqI+BYkZ2a8Pq8qDF0ofc6
DaZzkuh22M66bpeUY7NfOwGYF11IBhNxEcZBDWsmAoJPI8wuKDWmsUEVA/YIkNPzsZNejWLiCre2
RV5UVLpeeeJdLQeb/lphby1LsJlf87W8nUGxi3zv5US3VSWqhlNhG9XTm6PcfgIDw5oRGSJtp4tu
0Jnn6qmek5PiwCpxpjnKLiExQ4+05N5MMVdRs+KY7FGA+yV3oTFBWWK69kwskmQm/GAhbOiEYLSX
c9hTJFUDL4tA0ak9Wydzt9QKmGn2cMQbVv3VJJghKcjIKXOF+9JpijFpOLr4Xz/81v/6bUBDppYH
lgh4/z++0GfLONm6icPgLc3zwubnCh0iCnibm7xh4cfymHB7N99G5OFq85pHNfdh6orWB2kzEw/S
6OXvLVvC3mvqW9hAbN6ZGYA352EBRi1fFoO2fnYbqSPkMHx6Fdy+66kT8tDozkVV3L1PBjXNjORe
cvO8xRw2S5NnV4B9W1mQxHi6Cpp9amm58i4t4qSlxUzHiG5XFxV/dGjdUN3sEF5+GdXKbxCNmkhY
OnMZDjRNBshlkEwggLjWujHYofrLxgzMycvw0lyTh2yR5u3IVumcHY6i5/4LXYQMsm9gvY1eZtA2
xCBwNDyfHsaLcd+YFAftIjIWQscjcvPqgc5rHX4aM1mUkGsRCpfVPLFoxQN6DtsAg56a6f1k/IIY
OkMdc0Bb414VGweGFTp6qnSRbcZ0inYfI2AiuRpUONm4Mc+iG0Cxu2bcdVC7h10BetjhwehSXCgH
Q0Zv3+vZjfJ+UsKpNdAuQNbDjgnbJAiG9/7B9QDg2DPmvXKl36KDWrpexPU4LIRD6NqEEBLf8LV0
rnKpTjwCvtw+0ty1YXw941DhoQnmFNgO8DU0AR/57cDkH/ONoUmRavXnZCPdfFmZlIoJPqqQv388
Uy9HfgR/j5OcUALT0+5/yWS3+D5cN17+00n7O1hxntbqqa+fyGrlykbI59iDXBYq19IMNXYgOA6w
Q7ydDAGo5SLExazGb353ZLOO0Ht4xQ74yuL750C6n1luJ2ot23GOeqwPldVhUnILhn8OcTSeUdI4
TiWZyZafakF4WJtCaL5lQvThcVWGwAsNDXfP7caij1tJBdGh7kyG3sntjB4goWTcxH2IXWH4wq/2
FulTSN0Q1DqdU62Y4g/fYUlwAsRb6TRZBQg7Yp1da6uWJz8UCElZjtkhBkfcFZmpHWaA1VVy1bQr
IRljSwCTQG7IL97JtSiPnLHi5vrPiCqjkWO9/QM6iZorVLuZgYE5qt2JgSIO8EXzNTAm/zjI2lZW
hfjQZmnKaKR9MpuFRB5HtMZdwBp8ENhVfxUwjpofulKlVXheQJutZM/Sxu6x2JB8Ts9xuTg4r4pa
YdA+2cKdqxrmagC7nC7+7gNMI5UPOeRh7zGEwG8Z7+6SuSN7dNninf4Y1eMWLRPX4yNVkPU0XniF
2R7VmuF8VtilnyA1I1M3Nv+oitb38D5OU5B8FyeteRVv0BfTtRQtULNton6gj4t53EU/a0zn9tVh
Qa3Bu0WxbvVpkOAcnkLrWQbt0zI7Hu4LcZMhbHS2w0KYuJpC/srUfscjJKF/+rFEd8GGudAv/Iky
mlrM+AxxkhR1wH/o9IdkVRrZi53iElRGy9hQTTQjs2g9wg1Y76gj7SBJCrtJoEI+JDNPQic/J5cR
TmhR21zccTLoz5eCojV1E7zpUruAbYsFH+7kAEFrMvCoAPkNLKPq4GWmCEou67KPMcvYDpsN2a5N
8gv4b85bL3uETEWiVTQPvZPnmWWpbNFSzsEdIv/T3tsZ9SjhT08i00VX85smANmucGp3qIHtdlYG
kaSTxqxYOwtnyWhAYfjRig4PTHR+8Nwm8qAO/TkbH7T5TrOwEj6DPPNyTBJqPBW1G4bRKBbvSsYv
l6Tu7yOKWeUeb24do1JwNlJZEoCbG/SqwDM4B8bCmk/jT74EuGojiO6DokoWH2SxJ/hBPUTSJ7TE
j/U4JfhvrojxRlj/TYJtC6z/RoTrF/7gZ5a7no3nrGJ79eJaLzYJKgQfxtuRSsraU7U8qi0bPjoF
2QowL588urdlvgnXHTceA36LRPHPqyFh3paOhHN2XL2YPWz5t+PQCBslxmmhMox+bYbYXA8fXdUz
RgR+BzEi7Cw3enJOWF/d1J7YOa8RbK9H4bhMdNKZqtAG1CUCx4VBqmlCldC73AjpElEu6nG8RxZ7
batVTZR2lH7e2Fy5Q1uzMV+QcK9zGnh6AWuP8pPX9FbJnsCLle4xN207/JPzuOWsXbhCrkAT0coX
V/PUwc7GLua0tHTeV98hnsqcGi+wK/pUFZgUxAQ9zSHxEUryYFsrs2T+0q21UrCShzvmOMky1OfJ
8oS5FrJXa9jzInXVaV8aYpr+VNATunJ9V1xdGVTyXO90xhv4PmEW+s1KhnpHsP063L+WhifFJo7h
A7F/x1EtNgVnXTEXOhi9Zp3kBM0/JqCF2mpylZXzwtDf8T3L9/894ZT9GPSkUyccTdNEjisaWb/D
vuEf1xVRD1P6017BEWDJdTr4iJuXBOMKjT4zKcj4xnxqbDN/kkr2u/cEL/XMbtEhG43k9dZeU0Y2
JUfBloZI+cTSiWvaeeeqf7uK1MQe1qb2/trqXiqvTUHzCVK9zovMrfost4b4VFkzjz2sIaBMkLax
IXFeIkU/wSRy9K5y5pDEDNFrYa+nzl82Fr5HNhqA63oWhRppTfgthwC9XaT5/SIxNeED67aIryA/
GoouNAGU6NyOQgJZNl2YqSmClL0cN06kS37MBdrJ3oi8mcU/6/D1xmT3x7ut2p99I1sX5NmCSeFo
KVuUb87uSWhVTS4Atu+MBawlDsY2OB4UqkY8EXuDkFuaBqcH+hAlheM+dnklhVInQDsqh+K6Dlq1
SaDMLNiXzwTdezZMUKdW61b0evfDwTbKUrlXBXiOUqGgRFWlTRs2iO4mLjqP8lnjSD30WAPMEHlG
CWN2RfFRXZX8J4gzdNUtLOM3p+3ImrralRtL9zV7ysGq12V6iTrbYdByPZc+SWIjYaePvw1VACR6
2Gr6KdTgc4LlrOl+6l/t6hWhPTStR7TU1skXIix/qPdWVbjBw6F1qGZolkCuTvovcQ32kqb6wzFz
Sdj+gO3Vu9YeuaAkiCSgq6AlBkA2N2N8ZBDDcJofyBE1c5lloqQ4qTp5aHPVZPGIaixEI6V7/0t9
BwW2HvGNiDOXZQBLCmV0x8LFjvqqvqaN9ryYS2oBiqo0ddwPPaPIktKkGyMBunnMcpPClDBxdyoM
ZFT04liL6hV29E+5YtAkXymAhNdeV13GE8MbQrgxuBy75NGIWHXgekMG/SW5r8e0vaRYS6Okiv1W
r3ONq/4MyKlI5ohDXXZ7tfLMy41yL43gGldqqgfXMh1HuVjyEJhc06WLKX1n8zc4A4xmYf/oAJDG
ixSM9eiPsy1G7oTgp+o64IDfsynKXbuoI8bJOZUAJcXjGOhDv3lqh4PJuZlz6+3GwtKAI9/EF218
EAl9Jvw3XYSO7+gKCm0E5F1J5Cq6ucQ9Abo/5vhmOKVonUobIS2ppky8vAkdBSgfA/+1UzkaJF2w
2TZiQzVUVoj+rgrzfBBO9nND4mD9I6plfreTa4swgbypj/eVn/+84SquEWHa9p35tkxMQIlbdPBz
T1I19HmaD5vrY15eGj9OdWKz05d1hkYQtngtXW3jE31IRyxknWUbrDyh0DkA72IKGPv3va6iG9cq
V0rKevcOtiM7IyiZbk9lktkuf1cFqmEhMg3kY2dJvuz99E+iMHUrDFM0gk2h0MRTDn3jGS4+6+sH
J9/3xP2SNhLEf0oXSoxcgCHCZOCcn4bwWf+0D72FQuhF6JJQzIFkZUiTJkg+x33W7OA7R+L5nHNX
k6f1WgntC6FsWgSDRjhlmcM9xIlT6yKpfNRB7ySQNy8d8JEkTcyZoyXAPut1MMWfer20+cktcgo7
yHTbxegvpYkdjQlTQXBEE6KAD/8IQUTb7d4whRHOtdxKtIT1aFw88XXedAfBldGRYcqHsXKh9NrD
/7mGoTwa6CQ5ITXkRvVXZUzUw/YOwkDPgpEsMpWCddmmS3ghH+pBLSXDRuNoKHJdj2wYAHGxKNT3
LBjnzUxMSIMeMP3gmNdjNNcS6OEjxxUmaClUPyj8FWEalUBIwmtH4WnOGgsr19UFiAliZqhBdZfh
+vnPGZ4yl54t2r3/EdW7WR5yhxxlrM+CO8Y9u7g49rAigMoELQjiYXWuGuKSemdfbiF2og3LjOhL
PlBj8731erS6CqVy15LO7WZapoH1dC4B8pKn0EmFrs4hzrgyKsiY7mqMiWvj9HtrLRtT12apwZeM
hkRpRCnqYMRFPr6cqGzVBJQO0n78NNy0XDlmOgrswxNSgeqcV8A+kNmT0G/T5omBnKDg+BozMopr
0dPxEQi5Gr1s+ssBZHB2hHSTMqHN/3xKsRAuS962qunrAs2xGW0FLpTbuBRHnVxFrHzdxDyv3i6/
jYRd4WwPeITgN5LN7MBkNSRoOw+f9MOGpoV4aLWfK4snx//vMd5xrJJSwMo8Kgzf1E9KeYWwrkeE
AxnT6K2BUvtaDU8UDSxz465uuAT6FwQdFseUk8xWlnMm9qcacsXCD0zoev8UlKinBJUt34FR3Tm+
XPx7KnnWLdh46Fq7Z44xeltVKsebrfmoz+X0I1hFIYIIUd1bpPIUG1EDU1yvcl1gTO+oVa9lB7Va
CfURaDPozPiop1taC1Ze2V+hUHoi2wmcqoCwFRgRohlVSjp+rGCZ/NXGw83PyjdFude9NDG8u0gD
Bpfh3dLAOc3vdcPwv7vexUQKX51n6hsJewh2VoadpeLNJjSvfFR0PXV8JtjVuOl8C7/zqPK4v/H8
Vfv/3f0v7mUbq/7iLCt2risjPvDu0WXhlpB+AY2guAiJlyjEGY21dKnOVbZ+yYT7GH0STqYupeTz
0uD/82ag8QuqN02UVEFZtS/Z+j2viSe0Y0NF3zK9q5cUqPnXIke2vUJs8OxrFQhIJ8qaAMvIjL+Q
ixRWgT2OFgnWHlpgqEE/BWyrwATZOT60zbdXAIPY759tFUKCGntttvsp4Ic5kQa8y+BCE5BZLNvB
vKE1hNqrqGA7D4yMIe5lzvSoepZ1hCyQQ/0+W/MYeDxcIxC2Z0G6XbDqaIvL02S82JQV6HLkb54W
h65ZRbVeLyCex9QY6MnEV4FMSpF7AoeJdIUmK//69xrYtG5NMKlt9/RcdOKkA0fhFutD/7X+VM87
4IitQJ6BiQT3EJbNcYaQGk0lAv13OBB3NEFuHOV3KQlEE2TMEzOUPvx0y2un2KOtQn1IczZuyTvO
j+o7NfwOlXo8B1y6iJhcL3gH1uAOB/Q7FDWq/9HviUbq88KgGopOlIIBOYgqXULBtYNZKFCx7x2L
lBFraiJ18qk6hoOy/VAGOslbImkUZPBddTZBMGQ2+Y3u1goupLJYM1Sj29tCmr1QPtbCFvek5yiN
B1JtPvH8Y/ZO6fbdzWrBjncJ+7jpNko1Y5E2aJvi1oJyRrVOv/6gOziL/OSnBqQxTX1TsXCTTHfR
0JX/XKsT7RwDZ1s0M+D12oAZ3SfBZsvvF8B/DaQF7KGMxfROcfi+JWqqGxlzOTynN2kY9J67NpTQ
BIXBgI71wZ5WBGkvMl9WpPQnuc1mfMzVv+cTuM/9fNqtmtMkKsQhltlyHPPKE3w7TWWKzVnhy19c
vwroIWUQ8eAeMURcV3dzy46iAsZBL+BmIi+n7awA39s+F68oEbqhyDJKUw9M/AXCGLQI+qOvVhCc
UY+G4WBco2Unz7B5WhwsiX3YOIHZbm/uUPU+xrRlhN2+WmIKmKtOAID/0CIr4QcwRp40VVxWXWkk
RwOsX4SCnY3qbbqTOuRZmECbqWv5/bAhwz7z5Ufd5XVGIiiaRtMXNkdgOTAP4hAyj+KonWvoGbl/
jmPg2eXqnKhLwvSnSM17zgvPYedEeoDQJnH8+9TM+EqJgOM94LZPffwuik/GpQUQXjzgqrAGuJMb
fmJzTlQdC3t469vR9RuWddPB+Y1kTmA051gfIMUgWOIGAG6oz19SvV5+I9kQX6jxtjff8HF7L2lJ
G37a2auoQHcNIJDDMc7cT5Lo8TLH9P7CVyFf8bndlVWz9he0qapF67QllwLtJomsrBh3NfIYu2xr
Uv7qasN+J4TlY2vVay0pwMj6TG2v/BmdMhi+SIYCGfNxZNqoLO/ChuhBCb5HJdpHEbIPZcNtXhOd
D2/1emENFUuO5AZ+Thn6QJyckZf55flnzNDAxtSrd207D1Fq0IHvpAEmeifaBBmeH5979k260vg9
ItQMHTufdQo/PRDUWD4qdL8DW1xVLYjSVxUlSfTo/h0rPqhNkvD7XtIuK5E90qDA7crYKwXbMM/W
GFqGDfJH4WMLwJ+wS8egl58Abd9GrWQnKPpu6qBO2hf8BzfLhgMIAe+OzO/SY4+guObIhKViZnVC
uniMQxewgwXVUm1Qxxu9SzaMzRm95KZs1ZX9M/awm3DY7ZJtAi3M8RAn7T0jctbGCVOOp9RFX5FX
rO/afbRQ5x4RDRifynTbQV2UE4ippvQWdiNgNtAFCBCLX5JXmK0+fQuwOZiNQdigebnVJ25iovoF
v7qqCMNbiSj4g3y4TznstkPDUzGO6MMgVk7m6YUzDp0MzKNZirumP6XUtY7leUGQKleHwTLur4Og
ae8SyOGRecC3AV0MHNLJ6UCmT5LeJip2ZAiCOEW0UXGzzjjY4sFtyBnJLOJDZuMerFoK2+1uslmv
TZtWDFGasm5ks/qcH8WVK1i5NILonzy1uVLwGSoBif/eRCmLpiWTZK/2qLd7QPjDoMh5iW2CBb25
/bSR5QClgeedIMILIWQDnTaBc/yad8rtwSCUE2yX5CpswkjsCZBncwvkviWqtsFgc2b+kCMZ/img
+6j9ZKMocFgoeCZpFV2wKTiZLKanaojEWGI3ik5C5nrSH2D5jIGsdqpx6URsKfFduBeJtGElZ9Gf
PZdAwgbQimoDPnfZk+lXmdFmJdpQIwJV8Xxc6+7QuTu02z5cge7CBX4TTaLg4aBteLxfVJlCOmPU
J/LSZawMHUMnHOK5cUl6WnGr/OPwVDMTmD4siOjAcZiNzZ4yCpMlD5ZEJzduaiolSAn0Fkij4utQ
r2M4c8Q8xrJvu1fLu4rpnXKfOG8QoI0+XcjWSsTDRuDWFbSTEOQH2KiuNCA+g+kyxCJOtqhLkjGE
YfAg+NyfAgxic7LuDKgOvIS+pu13dZhDtvRfF0fo+dyskR55MpXIXGcHPtBN8Ni1w7PWVAp4hlLa
xeMkcXdUWwaHZUswV+s59DrP1FZpnYFH9+tLmGveD0kb9obDk0hQ5Za+YOERP+7EQ7cr7fE7h4th
q9WF8JbcQIrExrYvLTLoja1F6F5q2kxbh1e1Koaq2qx3V/kYbc6f3mbHKQuT0Ihiu68tXPUiMT1F
qUM32Mo//7PRV5tYh4qMmAOAhmsaYJhJ01qMEPT8r3wrKUxQ4EJIiwG7sl6jpTFHawXZjOEZKPWU
VMPztnS8tYUAf6qS4DNwxJDJFg6+6esEb/zjJMCV/XSbX20JRpZIA2uhx+mwEZVJ4eZdBKcDlPd3
lUQ8udPor86v/Lrqr6cw3a+kG7wtAYrXOcLRpzwWhio24DHEv06dLKEy0S4F0z38PJmXcb0ZdO+0
yHL1ShGn9uyAz/WZ6LFHTSOWAiGwakCO70Q8tDyiH6XEf03Mo7GfYgQ3sdwMU7v6d76eI+etGSxv
REt/yLaWW3L2n99WOVphlVDAvrQLr44L1f2prZMmgUP4lZZ2TBjZiUb2bQuHT7gm2a4KRCG+JcCQ
iggnjE0W53Ua7Tn/4rPwa9z3PicvuOAoEBmW/0ylO3dflWlHZWa+Ye3Bo6As8Qjbby9MeW6+qmtr
tek4pVK2ZUjwc70Rksfk5+yke5xtVA0137YdV+DVqDXgBPjH0FeZB+2KjuME4aa2A/R9yrtgGNdZ
0lXbq5KCVutP7BcavyoL62xQky33PERvnAR2NevGOXztmE+5nLSzi1A27Fut44FynyMmrX0I08hG
jfmqtEx9BgD6ClqgP+BoZ6Jj34DchQym6Jh2QNa2Gx406P+lZKqd3plCskxVeaKAfsV7TvVLLaAK
Rn5UZx0TFa3hPuU9XpSIzFuSLHnCCuy03MTun21O482XHbgEnU0rcVN2t0rQUgZ1ll1gLbI6aQAF
NjshgVikyX7gCH432hHkV1Uctney24W7HwpsRZ3rzT5Fu5lWo/oX1i3U3cEODK6bSJuStfTwwzHo
MdY2nog7353TbS2asHtDI4Uv4V4YqV6bkupGrGxgioa6bUenLXdF1uCYuD9ZMoigbRRB8hquZJV8
6LrJYU2DHVhAC6oejMGL/QNwA55ZHEGHMW9jMtY4ReA79/mBLUPvZWA6TUaXax+ZCe2cS+qvrhqC
/wRPqUpShGXiTmF5+Iht0/FRfC45rzRgpLgIpOMvsiuwEqlJ9C5NMa8ewK2/n1Qn1HlIZ8a1FYe4
EolcyCyRVJEje+t02rs9bSysO7mfKO6c1djDFku0lqrz6mMDi6KPB9e2w1EU+xtQTSdF7YcMVDSa
d6KzLpUfPO2/crpqZzHAHt4mJbP6obzGqBN2J00SQj2g9svu8D2I29Kn9TE7gtigvP8WOIxD1T0z
D9IEWBd2VyhILy9YT5t5VSRj34iu043G9w36Lg9PmLB09slZxSyG/tKKRoEFkLd7B5cCJeAq6TMi
YVC4ObbzbMLmpmNBQqyHTlkCuOUGS5K8pzIbmcHiDE5FNEGylZ5hYC3Zm+xhT5M3H1HAMd01cq5k
mlUmI2srucJj1jFUYwlQgxvpfxgd5T/YRKv1pliDLj2/v6r6gmRZBAyXI1UIPeTTcmwm6tqjt2R5
wmAGDcK1llFbWTCXtvF+5S5Zj2BPUOWtVNfr/S8uARQpZecJhcaXkFVx6KiuVqfPba5eB6DpwNxW
vYIOD1M7u+qrfDMmx6iY0wc/A67EmC41Vx5EDI6idG1vH/3H8N3+RsZBZuUgI6Kkxd58OQGP24EN
IvzObNr65oezWP4n8kt2xLRKFbh/5JEKtGz6ga0ZIcqeQpfqMTA17LFcksqOxDdTA6zK/F4zLJBb
b/ugqoajUaMSdszD76YJ3Jatn2439Xnqph7PlxN8BSJd6+ciNDCPzs1qZuUdur+3RsoHypiMMrRw
+fNzt5pYnCzZ6FdCNthz0UhPcEb6fMIJcqntbtTlkK8ETUsVD0wqRibbFESIQNRR1JWyq6ju3Ckj
Z7wNesOQHT4cJZM48IsN9A/PYaUaQSCjDWbcjzwL38N1zlQ6UNhOXuLYw5lm55oFUCowgIaz8nfy
wMegQ3yGenOTKvmQ1QMXcl99GneZofgncXgRzk/zakyDTjtjMM2WRTyLeHf418eYqK7XXXU1MC1f
+tfTOuVk7P/8os+o1vp31EvGBP2imdQ43/GLxgYL48o5fRTrub3GX0NlHfvZKYf9WYIe7Rvrmz2E
vFvePLPvvz3DeDVUvbG5txM6ysYlUpRQwqqNqO0HdClqBTUmZgOsK22zeMoSvwV1NpedjgbvM/H7
QkVT9C7n0sYR0V8aw4q7hHNlCscg692x7IHSHVKYU47+2/kQR6vpxnUA+xXgvD8ansZUzeLg7O+S
vVSBEQCwVVkreuBrIA0kL2eE6GkxVbhGTsjucYdYemnVz8wKZsVthSe30kwRzixX7VtrHntgb00C
v7Z9I+5sxYgqVznXcfnGPWcyPSGLdlEjNnmuhD9HAOsAsTnd7mKC7D1igIQPQdkwoQfhxmEaRL33
Z4GAWnzRF+eUV23GcmYvlaT269s8E03ybPSY6NmOKS2GC3/TASQsnOYX9re6GxEPe5B5sR+0f9am
50F97yXEf5GWBMnJDr/AzvtKere+kOhCPQLKS2fjTpTRjbwYYka1m9myWe+NidfSRiAP5Mdz0nL5
WBrGaTwmVK2LkttdKhRNfUR9FjRo8vWrfJl4V4QsP4nQ4XS8RVJ6+1g9Wa5b/bexiMZwK42l+SkW
S7FgLXJUFS5WJKIBRDnBgxnuLSS1yrdVH0NKPyo9qH8lGjxw8ahT8mZ63sqwgRsrTHIrIT/T4JAg
IwRhdO/w29ISpLuT9ABYt58AEhz20GKKe/tp++YKWqhX2VcjPLA6WonTPFvehe20VLw4bsTpF8ra
urD42E6YzIQQ7yj7QkZqhx90RfJHgZg7DY2ZcUrI26d83j0tWOXloCnucZgPnJywyn+kZBuSZvRf
2GLFDPHjEu8Mqu1tEewt5GtFV6B/E3XST/eliQcp2fNZLc7uPwTYheGMXhBA/mJBgFPD5jLghzNp
mtqwqvvidcEjwljwKbre4GCISxMooBKpMXzeBEVOronqep/VKVoHNDBP/jmvZn2uN048IPx2dAg/
e7Es7+QGIKeR9NvXtg1rDI2837TMearuGHQ3d4CAqqHXSyRhB3agB/gTSrDUj2MY2fQV3cRo2O7L
NWZpk41amtr2MegLcZNVnONy/GeXaSbALK9YPi7s20wi0lG7OWIV5FN15mzncBCc9YUh+JBm97US
eiOMNJwnntlapQ+9hFa+N945BntVr8KRjwqFO7PVudjsjcHP+itY6J1X7TzO7H6G37C1PPk1jsRL
hvrBub3md7dF/0RSAUa8r/8ZmsFS8Q2SNmxU/bZjSbbiGZ16n3CYr5wPC+9SWZlkAsCPDHFenAHq
6YDje5cu6iG5LiSS/M4kx1oCsFqXoHXZ/eTJMnOJPyshWw7meOsqPhoelZZTHzFapPKrzdQvQUWg
neGfFPSTiczyLEV44Ifd5j6WLVV5bbfgC1ZGC4tdNG031C5VqyyhabyO2fbvbxka+nyFz14tS93T
b2/GMrPJSvNy1G2QSBu0nPIfQaBOC5wkJvHN3hBBQbcTY76a2UmZBnl2r41O9cMAKUY9Yue/GA1A
wJ9ReREWRxFOJL2BRUysobhCfV9/cNpuXQ0ikB+qVC1/T1YKNXvZu8aKpJ1Uj0+W/bUFiendw0i7
vA0SizITArRyN82JzhOA7qP/io3EgUWDB/iXpnu9eyIfnX1I+qjyVYH9Auvg5B2XvCtb3E/YYrUF
GcCsIRaO9fwFi66BP5q+9ovROzK2hExd5d4lyNsADcHQux78ER1meIXIWyqaS0Rkz/QM9f3zAgnj
jg+vXewHrifIEAD89NML0ZOPNDDjkgn2TDwINzGHZS6/Bf7Ouu8+5VjxFBubyfpP2Rb3u35rEaWS
ghsjrcjufOEhDDC73UmifCrLytdnIwzTtLzCX/h6I8MjcnPHoZtGckhoSbzESKkhD8WEJk8+KHdU
rPDQEHaAVJLvBNwORrJUKA3SbhwAD/e45fiiLQHKqmEzEP7mXvxejrcdXth+WXuQNNTDaCCGpQhS
Wip6dCDsxn+96b22xaPEoX17J3E9nYor9kWXfc4HDU9smR4eTZr33krynAd7Bzox87FquB7TJ+Jn
gBcjngTzk7iwqGf6eFp0fXnUSD/S4YMZQZIfQvo/8FV1QcPews+fzrBdITxbbUEIVPENnSU5YAjz
PShLaZwOBP4pgC1+YBiBwHXnW0Wi1Yjk7WpagAkP/Y2vedGEuaWsZNI0j8fRLAS6eubEgnJ1bxQo
/O0JS5/6riQ5atDU0Z8jJHNDIaYee2YLrEYq40+k3GEr2Nez8SnbOJUKJFV0wuymB6LTjvaj1g+X
xaiBb6yrxvCa6+MdAvRBEpUjJ+534Ud4WPqbvXK9TCWNhNY8fVRAGAU92wMP7USzg43IlQynf8io
WQhNN5Rm9sXTAvWAtzz92UsRMWvAoMm9JB/SxAJWXCKKMcCnbzq8yg60XfHBnvY4etuipG/e/YuU
nK/YJNG7IekGmCTSdW5V5Q5z8k6fBS5OTU4rd313OmtgNotgTHVBuM6tkkO9D9lEY5TSr5/eFvrT
GSf+KoytPfEnmw0Xrwbm9lmusSK3xFcscsJtw7wuqkn2l2XrQVW23UN2cECAf0+R32YgT4kIcZji
FDiFoQq3GTJsXD4cDbG/DCB33NhYyy1KGZnEDmnxs2HkdPmGjdZ0FjdjYeMNXMQj/skM/QE6HMBD
o0bhCL+uXo2HaIibSb2lLAArUaYAYtzt+sLzOn8qBWNjMq3JtpquqKT3G4tBLPM1specUJSB51as
evAS02fxrC/kEL06dCiTN4E+FPAsILVGlxAPS/Fv5bGhkB4iTiXXRQ91q32INJ2vCkWPAfWoD8NS
PgFMf6qYk0xZ4q5oIxd+2qszHCXZviTeqhPNzCXyx5p02556k3IU2UQ1eET16gQQt3SeKD4qRgz1
87ZvnflIVgxTBknJ86IB4KVlkBnvtbZuBh0FLcFgFUPch6V6GGyt55p3LM14Jy/n8iX6WKRQILn6
GUsdOEBKof2N6aWzmN/ND+LAAHw/fQNhIUJjDqyRVQwHQdBn8HhkvRs/iswCuyH6hQ9yzu2RKpM3
MsRDld/DF1VC/I5l28ztr2cL2ZVJ+n/blQCx0022xuFH/DDXdcuPchjJAtSDK4QoGZHrqQXAlhvh
qpllUeOjxaVQ6UJ1EtRTpqEoDoKRi6LZIVWUP3c0xretn1IzDvYkvy20t9CP1I6Sp85UWPTkWGDq
2pRCYNmovVfsaViai2nzUoWS8xu6/+Puk31jnr4y1bvthG/tEJn9kSeRml7R6qGsvAaMeVI7CtEy
jW3wK9tdpK2G60SW1tHfzeTjouTMcRhO5t+WE8T1lTWurGvVNkH08/t3FsC0j9pZtjoPUirYqpeP
OS0VIOGWJD7InAVvBfyw1/QOL5I8c9UXvofUL5opb7R1UAQsdApBf98L2HOPUwqks6iQrBmLLWzr
Xe06yeyVThktcUK6yudoDnOIWNZkdEjP08jUmZgQ/QnT0ufr31NJuzim40DvjHNo7sA9F2keL5ie
A47QXhGfUyRxfNEHB0E9rDEv7hRmo8hlT/rbyX1jEI9rx38/BBiJtmX9ABw5aEugQWbSfKa3e7OB
0iTdtwcp/lh5loqSqMVXd7DAKLz9HeAQjg6abd/enoBqCQCkwZg/X7ui2PT5TJP3z5HisrbjYrMB
XQdruCEMHwZvqZRo2UwN3JS4Eabn9UYHSkuJNYa9zeTa4H7TzmsFPv+Yt2rLFao/MPytCZeVBg1c
W803wAHZFLq5hl7TYVquxWDrWsyPpjELmim/JpQvzATSDNv+FPLO165GOwfAT/xqo1Y1vrWFAiBA
Q9ctoJNNmYqjrRCmvi7rxUVPAPid8m6Ub+zQA2KDkxPGAkPQ59NxqXOpvE3+lpMw9gfT3t7Tx0sK
WmCVCUGvEzMmwGbpIgVXSHyKmhwBzrVmtOPGgqdSQIePsse8Qk6YMBr42eHoysEqyMzMkfJNCdId
YMgj8SXjCfUfkanTkPwhUpvnQZARsDF0hLzZaqkShogtjbdYlaG9x72XAxnRj+IavMMEXs1ZvoT3
cS68DHXn/BdgPLDMLmdipBtibTSubICNJTRJkCrKf54k+T9jqWWGza8nms83LkiQKEL8qxlqBj00
T4am79i6gV49ebCKRCJrbtrtJLbRAOKQjHkxm3JvxEZolW51towx5G3Luzwzk+AXe2PDyFfLhP3w
Sl8iBGqB6aj1FAo1o6eXpHV8C/XBKhHjF95k/3DzERqLpht7cFoFK0AtFV1cyHxZp/Toc8jmvSuB
lOMyXMcfNn5omSSvPLVolWyzfDO2jrXyUhoTmEfULc4XMLqv5oSNTj/7JDyrGXK5WavDuNne6tMY
1gff/bnRSQ/B00OLfB7kYCzxzSJ5SdDt+Y47tjzUhd9bjNz1icEQVsqXiv7s20UIesMuD9Hdz1LI
ZDeXJjJHMeHEWVmKrTqqL6/r89iSBcwCDB8TKQcV+uGHfg4bF+2R6Y4SHpPaJYLMdc4xC9OfWob9
ZvkFVq+d9ot77p3yMRg+AUPqhoPhWCPn/b6Lm4KipgLbIlXfq33MtFtuk+eegeGuAnNt2mPvjeAk
0YyEgxkVBKfQD937u9/7aaWJSougVTj5CHPsGpHWbxXhPV9A9FbQXuAdnHaqT/WSvLCrcua/oG+M
nzVGTwsHYF4xQHEr+hwoSqyO+kE7b7d4IGF1QIZXs0nFOAo164kibA3nMS89VwzJMEQy6ROtZiU0
ZHjYFRvXYYjB1ZF81c74KEEDonJQLrtdkeQwc50MSDfG+9e4POwZIjSkyeCI+4DdwPKZP27K/Hr4
CSdi8r5c1TlIti6jwBzO9ripojwiTq5WteK2Gx/aBrNq9iF9e8GgcuLykL05vSWg5bbzCq+rkMSZ
IryKt2lTWwJ42JaG58Ng4te0HY32lAjhRLA0Gv4hHX4gsPvOa8WfpG5E7KyLF+xpV3aR9nvRTVPG
GD/h6osAI62xVI+TTHLNJTpPG3VMlyvPZkjAltSL2xADBTtpSmmgzIRCPWdg/N08fzmRzkSwWIGm
xxUMTujsHJBHVpISRWRZARjbKRb79yHC/pGLu2EQCLMasINnQ8nNdfwpD8Amyjb1hnG7le9Y8rQ9
hxYcCKtAD7Z9e0mADGtXEysIYAaYVYat6ctH8Bd5nfX1IV9+hT7BO7mNl97EmrtBbMJeL6Fxqmna
xAh7PNqNuuxXPSl8IYDOfUGYCZbAxqcu6CWmGHvsB7K0DU1TpOR34HyC2HrlGvm5Eur/aqwSGSgZ
b9D9Aozx01OF9zBP6RevLv2Zxv6FC9z8KT6gBUn8pH0fsNBvrUX7CgekZ99gBHiaGFyidyqn/8st
T5tx2dgv3UjPzLfrTkjQL9N/8YRQIcCQIucnfWmvTHxad3Qf67G1+tckI5VfgJMjVYfs0hoO/YOr
Q3bzAXZKnTIpTfw/Edg4MDM8kzrS4wgeeWkj82ojJkEWuFPquvnQdR6UtM8yR4ap9PNx31ypbm99
CT9YIjb6lVBmIMMubJJTDD+HHhgupqhPD6YvT7jUBrWRSIVX4045H79xb0p3LqMoUYANtF3eKFFM
aFMzG2QN0o+ZcxvHSYyl2PEwkbWLF90kOZ6gpkMBsm4kANv7Xk0b7a0V1X2BmZMHbJT2l7r/ivPZ
4LtwJP6Z+1FtVBkgeck9KW9JpnK8ARW9CWYfn0TOCYNOiKDO7/dzjaz+FNFsqKv1Py3279yvOydc
j97+WcxS2Lz8ZVa62Wc/SsgvKUK8fvMJS0MaGvC1c3bARNyQH3oAmOjVzQ/LgtyiI5NbY5dXbsFk
fxIqwCnVXuPge4p3CSbfsQRD99x2UNLcTveuTWqANG0wENYW5KRzDP4LrUkghJt3stQ+WlP7DuWi
1JFwzU/4dW+EJMBJAHKrPYfkrKvcF3PBg9Ep4dWcByijawoaooVU11v9wezBE97gOmccZ6+A11jM
zAbxw11tRSCFJfN5NIYhGtCWHxArQj/3NgTYhBCUKqIVz6ONYcaxLIR5FX7/bdz6lcdj21U6A7uy
QpXW0cRmnviE/akDGYXjqBKoZwMdGVXKIDOyjb0uwWU+7o1u9+bvP2MCCbf6tycCBDJIDhFAd9zM
kvFEoLCUo2TXAcO/rI3VYbtIdK8TLEMM1tiSA0NMswDG99Sgvp9RAufW2t+uY9JN6ZhsNQEezoDo
KVbvIGSXJIiP037s5F8m0V+zEZPozT5X9k+EaGJDZP5UV4mbgBResEZjgxU7HYPiQhzqF8nlDMZC
F8o0gCZ5JMblvn52WbLYv2oqrCbczl62Ase53SeEFzUVE4zJGWMGEmYlXb3UuY1ngKevZ5dbXVsR
eTpgLhzlXuJTzwjGodThbKAvcvpiLNj6g7EfY/MjqtrPliNj48Pmsgyt2ICaBRLOhyb0qUSTo/sU
He2iRPAFtpnHRAk6t19bleck2m65EcnWWFgB6UiVz/xVxtxPqTMosWroiKHOIrvqVImssTxFRI7Z
+vv1lLKSmSKqKi+0CczpONa41jRbGYxIpPUCap9u5sSXpmHKqnihUp9C9x3eTU0XoUvt9vudk5oS
RKyD9pPKhB5rneNZkuW5VRXVSe3SxeiqBmDxGBYG1xZPrGH8/CgSVBZHgNArzAJfEf8e8zqwwWr+
u1PmmfIqVNyWR4JBwxzrl2s++UX54/Qv6h3aRh+8tPleHezTxvw3l2Aci7m7UV7KdCdxyxhE3jPV
zqFVsFBd865NQJnbT6Otdq0Ey6mYnReqadGyEYXUmw+LDru1QMCHV82xKmxsdD0CfUYKLW2jWgIl
Vw6fhvUdSeBm9Hrb960NDCnIxaU83NjmpeXP7uw6e4AbX7DmpEmtk5lA+sSUH4e+ECAbFcoRvuQ0
5lT9iTWWx7amAls7fmsZzGjfuyvKkBOkbyGuXGGLLB/QjHvwmANXoHDqtsRWz73yxWjYPjAQjUcV
x6Z+iavZJuaxxMhYUC2WGjzFgcGpAyL8tgXiS2tXemPXIMuvaUAcfb85usJe82CKG6UbXFm/Mb44
U/r9ixxQJrIajA/u56CkyPzkdisVA0Hnjlb+U14UFAGYp7yNcqQYSyHG+tI37pPFvRJu1Hury5qv
4nkhFtVPUwdIeOCeaw8n47Bd9oIqfBAWX8yenYGUPoKn1RLODwk79LFCQyLQmFwXuSCSe42KmBUt
cDaY8ayGT94yLKOVVVa2LtsZeWJx1AbzZ3jMb8FE7f77uOegugINHPok8pLa+rmDN2W8AaGEfW9k
TPDW7mjnMyQTvL2W6b+v8t89cDDaNh8wSzkF8lRNQb24/Kp03qc0J4noWpGelABEJitHcz3KNhSs
77dGloSBdQPzDSrfr9bnO5ijUISXrprbRTJ2GIOEnglZGkdJbpxZqwywY1yfuIlT6CCRfJZX0Jcp
TyghKa0ShVmEmtosQXXb+C6nNNC7p0Xv/Ed0GrehyG845cfaqCXLYsR/xzRbcp99DPFkQBi99qyL
n5QYey8Nn7lq0iGVz6BPpkodzdMya6IQIwetOb4SAaOdvwO7hXwDpBlXkZbZ7s89WAblDuLXGScl
CRez+Nzb7WSzAv1a47DIzb/pqW714XVPfvQy7+4nzQL1ADpxNRwwmkWIBfSFHilxiaBhc6o6iYlc
T0bjzDqkWQAZh4XMgtHhgDcByHLtwLRWGyZ5vQP13VRG2bHCM/AOdyKGwTjyOUwiNauAJm1UZUka
0jhXFGlLES/otH09JBBYFywbogonF7BTCV9cSDxCBcrxqSRt/z83JqnnpDhPiFng6rHSyoI8ekPU
sSsT3o3HK9on4Q+/UpGXEQQmD/TDLk5k/7rb17/0rb6asYA+kBAcuqqAnktTRJazdCXHUHNItphK
Ul3nhftaaVXdONEidCEiacdV3SyDmmA3CfBa1KEB72OQWh1R9qzUuW9tgDj+TkHhJl+KBznP7ukR
TmLDTJOWo35+CyRoX2H12KUsMe3TDFK1/0ctf0ioAAh2CeBzZjMNLz3uY1S+iZ1L7nsGf/XpCx4d
UgeGXpE9ukHqAR3p/91rOvi899TKC2hB3K6lZaN3Ui7pFgbZ9L7BSyEOXHcDatYIb7N01SxjcKeV
8dxPCdgHOeVS/3t3Uh8/bQtHQ6/yEfztAPwlZlN+3waelN6YwlI3HlpOV2WwhmxZ9XTGaj56mu+T
RQ5sblRTYO1rl/OMB9zXQ4E8hy056d+6Flxd31wM5DGnruH2UJEqxWXrrkII61pou4z27sfOveqH
99nDDi9eNL2N+fIaNtBFjFcEi0D2oViC+ff+JkmvJDL7IXsv76XKRWxASKY3o9yx+G8SRNnED1oK
nyWRL1MEzFcG3Xn/ovGq2FWiueqP0ymw6eJSW1SquQeHSehCjk9xwiqu1FNUvkkaMZvJkVCGEaYZ
QPSxLRNhE46TGRz+boI4ZLRTo6Eu4YvpCTnyHVJyHdyesGA2ZFK/IXhjZQA0/rcpBU++uxlP9mW9
kUyDr5iHEMts1q4htPOE+y0gGdTSUJitbFJ/0BIG1wuFQTZnNjYVfa9qad87SR+BYIC7tU7eoKqJ
rtEuZJ+x8YzTctGA49f+FKdS/7+Omu4Okp38Cu25RIFOM4CxS/T43E7MS5BctDg7VvDdAIiu1+RT
fbS57yU8j5uLxasxtvKOPEuAcFCC9tzubGCgU8ScGhbbeGFDDJe0BBQQrBFgTgI9OrohzqmzeGOA
n8Dh/3WRmYhTIN3fcfP1Py+LyTXb49uoLNQyy7GxTUDuHmFnhNhGatnLeD5754wnujwICT5mzldA
IUncxdQJIELc+4IqAe10gD9Ifjt6mkV5pZxfDtMXzflB56PwUzoSTXOAwkDDnM6+8CGkrNAFaP2U
14OMmsmGQ4ZNEoK1K806t8P4KiamQsre50wxKqh44NfCdyAF0ohtlkNPHpooMi8U9dUuuceeXuRz
bw75cf8BQ/QGtNBqYQuBBBDx7fvU+gZXjxSjmlA/qoBAoDAukwr6gq88QVRJ8I4E/mPyZ5+OyZgh
ol9ytsLpPJ66TXTigtEHGzHXGtruGOgMbrFpfqVo1D+o0rCHSSTpBAfhrMdj2ujHpYtaFTkeQ9Kc
FXiCMIeUsS3afXzpqgP71PWvwkhuQgbzkID2w+orBwDnpNidVvAnoHqhjdq9f0q0qzaZFu9FpLwN
7QN1Y797s090sm9UeUGmiRtPSAs9Aay+bKlr33s/fz/0NgXp0hFLXRTt/J4uWmD6w/M2TMtgIcb8
wVIaaKHqB81tS2RHRr3wQc0DZWIOaXsHjD1H/YXgu30c14TIL70AjN5FFc9+aLcaYli4FSjh1G7r
/ZO50Rlx+FdeEj1RoU+ygryjJNZJZZQUnosmDGRZTOuYDPYw9a6wjZ9U2wMzt6pZcbIHferyeQOu
tiyv//IsIJ9HsMIflDY4vzIb2vCOePu8pv6IRp8IQedhJ92q+qV3CY7wqj3rQ13hDYvit2+1+13c
9J80A4AkrLrtOsHFNES4cLjagXQdFNB/HeFpATrc/kE6sv6irb7S9KwQrHYYfYzp5dg91EDjVtAE
FOu7jYrqEDdm1D3ruQyHmNV6CSEh4gblnBCp1L8+MwYAR+fEyich5CjOvoLiHH/LdxBWXdNMjb4N
6Tr4vhSWnkS0rAvPvJtNVJ1uuZ4UAR9UWi2jh+NlU2LR0XsIVIwSExh3gEqYhozeX7fXyFg0Etbh
R5+URsQQwxVzfaSB91ppIvcGwcgD0ldebY2bbYl8Oe64umcQAjSqPad61cw+9CH79ByuDbhkfKJV
nieFVIaNR2BvZ2Pg917peYvLPUDzcoqb4yhnp3w1YxdHjK7WnKOB8gxjAC8v3+hZRam+/3AJ9hrL
TNaYDuTp5Lmq43Gd4Wr4vtsuR3vu9qQab2h0QGDpbhTVY/0UC1PVytMycuyvcGgWual/TCLVV+lZ
kGFc8ZLWD2GJNOb5Pr+sYPPrrtEpClsUNcHcVDMvKWAF14DBI1E/5h24M6ftydXU1BTE+usiEwAf
HDkDOTSZjmPMAHPwOWJGxQ9lSO49JpcVM2EUVThf7RYcRUPcGhNYuvltECwFjMUjeDSW5VU+iEgy
2cAa4akbUW+9JJmWuibXA8IigDksF4RSY78jzc5uOUXnLSlsFAAODwsEOI7LGLGkDtOmaPRDvrZI
255SGIpjFcSsXm2uCj1/w+RgGIndw5BozlHugALnLv8ris7DU83ztOV8npZ+sAGWGHBzgWOW/Rx+
dND67nHFp3ARYxkNK97Ezgi2PdwjjVQbNAaSGAjCYSYfbeGLgyTH18AFVk1H9umI6ezHUgBVww+j
ex6q+yFduseF3GfaM3GzktmmUUQTWk/aHXFI37mv8nxY2D+44k9fqShTwA6Gruz8SJmoEG8uRA0S
3SiRtgi7x23HQe5fI8PlsHGFYwWcOOFXl8XKxJGFAv8ThvXXvmkQfqvB4KjtzViV4F1ut28DiK6n
CsV8BQ1xwiJhvbh8DUeywvqfXNPTcB4L3FGB9izeG/Ev6WJlUpAJHCJSwoG/9hp8X/w2I9iGpoOE
dBnJgY9YsUA70nSD6sWLI2tSQ5X3r2qsyeLxWZSGWY2LslovmQKovQSRLKLkjYEnnbwj3Gy2o4jH
02Pip59A8IbjibJ/dpcyuu7SWPtYL2rwOch3jhFJtwMF0vxykBSC2hW+TB2fwLLAJ6VPLfbEb4S2
3SdMUWae84Zpid8GFrd0lKodpiG+S5wusy3r2Nvkhrm71OzhSIo173810rhqyVz5t9+dyLEXNbSi
MLA2nHkPLUzQjCQVIjPkmIqSDZog1unjKdsjZejjIV3U05snEIurWPMvP3MATdyr7/tJPkECTe5c
7/X2f5wRlzEtlcZlGwN5K2a9f9gt5iY2MT+cXgBGDWobUVTYfNQ/MeK3xEY+rnBSkGOWSBBKXvuo
KTzsqElKs72U3QXMnFLXdJfABbFmUAaI9F0adLY739xJpHRTFjUQkwahdgLL1Fa75iXOeq36m0Zq
oeSno3zOF6M4okgfmL0P
`pragma protect end_protected
