// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
CJIbPeUMprDWkgPHC/xWsoN4g6dUvtOaUdDRWkLbjOrsuFzdfcNV6hgLkn0GLqlX8IAgSOwDpsLy
EIeSjCeGYJ7bdF0Xk+LDGRL602cvtwY++8HOfAUjZ8+nrOel0I+2uEGz6RgsMH2sAkypEpC+6nz0
Rb/M50sb4j7ZrB33c5USziv+XTKVbzyl/IzwVEmjVVoSaQW6ST1J+H5ugFgC42WmQpcFp96F5Ddg
yTzEb4Fz/0BPyOeNlLXec2jxhnACdMXhqd9GAlXu1MmO7HcTHkYn2QZxzuOOGQa1f7+JKbOKXDUq
9+43u9nth2c+9wqOPi8kKBmqHA7AvPEMx13ekg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 17904)
fkFNrEdyPcLmVqXZmCtZ3wMdOebi5c4rbL2aEk5IUomdn+pYsVIlVRxwU2GHQD89q9JWsq8VXMgO
kGm7PhDWtvjWxkDH+OhXK4mqB5kFdH8bmqsRFQITX1l+HW6DoqoLLzZQ3t82cWwMJnTLMFVj1v7V
ORqOM+3/JfmCarQIoALXbo+bRm7Kq3T5FDvbTnWV9iWmS2FON6MrNFmknFgO4rYOTPnDIKMLMQ0X
qfYDQ27ZBzkniBe5EgLBcXQOe1vo2Uoz7x2HuD+rQ0dmBOP1UaxZCp9oNAJDomIBwN1ZPXIiMqAG
Cc6NxNLKgINYpabuSY2y4xCCataNvbyi7LL23uFsqq0UnTQ2KVpOIEBZK52SXx83qXJgY7ewDscB
+EwKxnduE8Dww6cP/iMDcDxwbgmCL3c2jS+1XtYoAv2oq29GbNRBh+n67w200QcvFVe065y42FuS
xgQI7ohbfbB1B9O/qbVKFggvJTIO+kCN24oQyxzvELvchBlrQ8iWYVIhPuieStYQ+XZdjL+Auo4J
mEN6v8nP7Uo2w07OV+f3gTG6ftPO19f5bWqkzZjivTF65a8tb9cSDh07fsczzcW4EdMLHL1tdSwo
Z+O1XfT8NL2jvfmWEXtv3o7zBy4oQ6jW/ZA+kN6gZwIk3SLzE86pFT+C2BQoSnq7GQ1PP99JfImk
04vW/JFkujIyrCptv1LU6D0QsCIuCHgL9Xf4w870cSGy9/zKNnR+A9iuyWpi3rF83EOnKyX8xoXM
4FXfzxOAmc0jj+q5C2IVoJGvX5DLSSKnkhZSzFFZNcBEdyH1jCt1S20+CflMi1rfbIk4q8nntvum
9eOj+ZaqaCkKJhX8P+D63o+jB5i0boXp0yAGH9EKgSth3T33nomQkhEeJzSG5ihkqtzOVcyc/YN1
tZc13xCHBbr/haST1+5G1Jb+/j4VzAcakO18vLCZlcITU1k0Ef+/N1tvquaN22TdEq9zOEOEY5wO
cGGdtzGRlSOAkouwuC/TQk1fOc8t8XWv/6h0aOXH7kXydh9Ej/w3B9rznr29PyS8kw9QQm5ALIDR
JVFHsg+JvUQKf2PB7Wu9n9YRTHJYbhw2J6TFZwZtpjQJxpg5Zi16g14eR5gw7S8p7IJ7d27ByaTM
mYznaXxjxdIIhzBh2qJkWfSut2VTUeTV8LuWVYwLIBgkhRDy7d8ECALPMHgHVwUCo09iowWfGRaL
fRbsMdlg2geiYXa2w8kgGyd6xdJYseQg0eA4jpn6fuR5jW1ajDUG3NBOUHmeVoLcRhIhzaUbmWbH
2ljHBVivNdcxD18boQs5P6nnvm20I8mEkNfj0a7CbvligdGfdoyDFzQSAnU7aY9/CZRN/Yt13lM+
+ySxUOQ/YDppIg8VoKinIvS1CtrH2AgDW9Boy3l58ozS6I/x4u/A+0vwORB06gh0WEHCnk72+kWT
6YVDDOX7RhamL8hLJ8Fr5Ow5oCsmYK90/LCwpSknjtct9OJhrcBtCpNsM8klb2xVD8IXOaP4cqKl
tkurKBXtJZn0nvqJT67vUaTYQbXLzdKoaihtQrFVT2PvmzYoZdCiAsvpnOFmeJ0M4c6/fqKoEQe/
HgxwYFqAeIbhD7h3FS6ZCezEZt7EnJy0yJBuCqrRv5rvPm/N3BjyQdiaXT7r337XsHbLM4Qsay0m
ABKrxJZwIkypJmN7hGdrHPMihMWcVFmzlCfJr+yonU6M95A0BIrtJLjaI2U6ccr42ie+8ZBXfNhk
/ulPcF9Q2KJIUzG9vjb0VUC3vKuXMfpB/ENpGJkke29hu94OhXt6n9vkDa8HX78jTlBFNbRREx/L
FazQ6Q7cRLHfpI+s9UWDilGjrcVKQ+DZ4aS24OQxwSeDpthnecGyCo498Ym9G0fir64vBTVWp/xO
kevHkQMKFDo8ypdCaTomlH7nbsyz1d6OnYP6+NgG5EvuY/p6gds/eaq8QOUnoKN5l03WA951O041
5AoagvQ2I63m+Q9Ta2WQMKdglp2yUCkiQpJMKLIn6khshGgB2gQCFLC3LdtO7WEDZMZHMI8C+g2h
H9Co8dmN6KDsNAj/pimlhbPLAcUcK+VPMgv9Y7/uuIAfvCL05nU7XWh2585lh48o0z6UacW3IL6k
XZbNZetGDB0eFMIvIVyFFXk8iERa8uAkIPVzRwGVxaxtHAxPOFM2rGpghI8bbyQrcMUQYN9U2ZNg
PtxfQEtoNhQj9OXgO7gsxBLa+u+MiWD6eYnj7O0J+o0wBhVw2A8gsaScKE+dfj3U3/oL9SkRPpUq
6mVctBybVBn1jSTHGyKykkFQVq6zE9iX7X958wmWvQBb9HJnVi2nd+3WJI7eKbauj964KWBa0w6X
ixB0BjXyPEOJSylVA87c15KGdqI08p9IW9Gp3+R/7SgIy/7xH/dDrlXE8h1uzZoZV0ABTqwfYRm3
IoiQ58IK0/sIqnvBhuT5RnL9G7G31GRKC2gVDMx5Hqd3CrDOMr2dCt+Vs0k/tr5a2yI/aX+u+eTl
K7BBVb3LjYsTJwAbwCEobesauLWZg8FkZT0rwXKaa2qJjm6zbYCi8RfzifKZlzcvpXVMR3X/Wate
s0XdSoH3NhKIOlGlMFQd118JuGBkbqCT9sPBPMxc5RXa/ubfvyFWwrZfHdgpDlRPiiids4gOOac8
i/nB3NkT3SfDobikTX7OWzPdZ+6r3spJFQdTYEMjivg8J2Hg3K+DxJV8sJzO8vKmLOYj3h3WGiwz
BJwhSdDIDFcGtWQINZaJ4w7vru3F9omuCSLfxgFXYtwxFkVfj3nPZPh2EU97BREo7fQNQCFhTUtz
RCzk0vUmnJdqxwXqzzdaPaXm39z4w5NfG42TAxPIyzl3C4f3E3tYnKOWvSPHTehmz0VJ5zLZh09f
z7phrLE/Jo1VxujSuQkbQG184zQ82V/f+Rnd42cw168Np9HpnUDTmKhss3qMNrEJ/9gD8WxVSO2e
Cyuo4kqlUxbm7Fl2yL47kukInZNq8wPYN+IcjVKUhT6PXr71H/Q+TpEJUPjyYRxsNkdSc44epX6S
Qumh842UruMeqWfTgWI0Aj3YO0pKmrVU8Cm7RarUyXDUqjKAl3++lU8dlDjt80Ac3AFtIXNWEFtg
ZIw41OYPm6AKbvXEJHIBAFZNDc6i1wqFPzRTqjqzzeVN5SzLZmno+RHbLIZkGGzECVCYPEgilUDF
4diJC55dXdnGEdJhNhe7Rg+goTQRxAt1YcjYjctB+D1E3/3HHIboltWQ9E3Wj1pLMzdqEFLjjerL
DemH+Tk2SRAGwUU2PPgyWurRMzGSGWmA285KscRxkoOQT6bKddhVdcR1hB4y0NsuHV7VMHosGyIB
SYfNjgh/A5P4Oc5BrcHc6dZD4B7C3jEk1Z8g4JBjIG4jCePbSjUZBFd0Si4lF6Wz7Esnv0ibJfz1
DmC1KH7z2i39Bm5RcrtrxF73YCY0nljoHiyxpryQisyigv9C8dLMMVcdpDSsiTrT3apDToLGaB5A
RYxO4yStTBwUSSzP5cF5qSyenEKAkstw7aOCH8e2pquS7ATMkKPtBPRY7SWg+TCWA+bxHtXcoAOz
M4OMNpPD/fQC9NZ7mZ71LlrkgA1qeX5ZKhlHFEMvhse77PjBTPUA+dmGZkbP/GDxLLndC4nLLGkp
zF+gc6+4E0Ny2bv5fX/eAS3uaBOWb1e6G+Sik0t0UoJZzs8tQ9c1KxqPOpNNSll7S5qMdOnWE3ea
drHewktAGcP8vBIcU++1rvwCNa84KBe4SbCrThgdddPcIfUfMFaz5LJd0KYQlNbZ9mMSOKoKWYrv
BLEAeZfYGxSCNHGf33OmAAzZeIwCN5g8OT/WHSLDh3UWAnH+GsN3kRhFa3fBH5GLEIl+2TZe7hI1
r/inb6gkSX2+fdt1APMOAjMSP4EwZ2RVraFxR2ajvRi6Xx5cCH0VvrPyEc+374oGmFoXswrS5YoD
gI6BJjWflu0egE1OCJp5d3acoex0A9isMsiB/XtJZ0gtk9H6B5wOZ/ZFjizv9u0+P3z5Z94KAsQh
6BLI/QtVmPlbxKNcWv+kwCnaJLIlw0bKoX9yAI7mAKAomwfvL6KFjJOF6VqAeo3Llw4VLo5fqOit
u4NZnenGCVTH2YCsWHf4rbeDsAGZxcjhF4mru93h9PDjZzxUaI6N2gIjWkMn38NWi4SQIiH8qYld
z9jzCTx7FXql5jAlA5BdDaSzqzqu/6KI8yeDngaTA/Hl4aCdgUz0VlPsMcqlYN8eOv+4Yj0PY8dr
OOW7DAhfmIckaoOAczEyYwE0S26H+tY15LsQgGKVyBZnUQHJwe63UhKFLtrDl5DnK7PbX07J40Gi
h9O7wqsX0Ba3xPQgQHI5uOsKCfuCvm2/EzmDjUWW/Rl72AtwRZRGozw5O5Lj4aLlkAa9hIlG19yK
afwNHYlwXKU14FufrABCrRueGGqaec4ksFDTOK3cOwZw/jYmtwkIkmltRMapg1WqdTmqBn+xoUkM
2Fx4k96a+KEQyBTmXUrb6aQkgSrybeWZqszDQlH4IvqBvaikHq9g/PFr6IWpdiHveD+I2CFNGuPr
5BaTiyPriN1lE77xNeCt/qy9BEJjb+MnHm+nVbJAaBjwNFSEsTF44Key9qZqm+1Be+McMA2o3h3F
iW83U5UWbQxKqAttMkcz3PPlJZfuqzGbhO/LrfvVO9BKvv+M7Dn2vmM45TeRqDJkEbfsZPAelv8/
1Vwtqn9Q2F4VqW56Ae/ZKHRVXhVtkIVPZQPYnwFnPLZIxWYlAMl0eN56Hj3VrTaz5PkB6FDWOvLF
0Gj72YEdDiZguTs9rNhabCoN1wmaivNi5wXWU2dJLMhgP3rACnTt1WCBVahN7QZWwHb83qDenqoh
ddBFMWDzgQEd81euNU3amyClQdWLtxg+goNoIcQJ1iIYhAm22aVoxCJftSz30ZZjD+QALy44ZlIh
UQBZse8pPos2b0AntiYarTdbHuZrI3/xyxV9FyosoAIcVuRASOvJlop0NIPXBWQNYYfyB1SgvY3D
4M1Lzdob7MEGtyj0zF0A5kwG2ey5EA+9Z7F1QjIBiYze0P+bsKazm/HdBjwWWpgce+Grs0WSgcDg
vaJXF3Hb+bdErEoRn1V7Ln5K12dat2kryWLOusWw+xKzmlx09Aat1Wb38RIPTVDiyp1YFoksatIc
jSp1l3YmDqiEf881S8M9xEs0HjB2fEcwpufRvdTnVJExxPVN1UJrDfE0TXmRmh543pTduqp/D2DW
1bspfXWXxu14e/AIwhHkruKO+D2cyY+Y/Ogz1WJhmdtXeNAUtaWcykZYwgFHfwtD1TnJqo+Li3Gn
i2a0ai0kFwj50e3JPCKtPoQFuXEug6VtZWi3GaXMmK+CnxAOzYM4iWZs3f6Ipwb81n6vyi1z2xBr
JOWrhLrEu74wG2BmcD3ihgfEGg6fP7irb0wIduIjSMRkmymJoih4ah+HxMW7n/JFfTq4qdbGVMTP
zcwxu1GW69hNtMpNQjl4hKbiEemHJAwYbUDn6p0ykU5wVmWRCSYhfIlVIRsFlN1JwWlRz2ZJgTbZ
UhPJOsnsvilPWC7UtoZiEbHJet7N13NwD4erkVLstnKmIGhKbgaBizQWi4k8T37PMqiapvCv6izm
OSyYA8+zJ2Gg/mYXkXj0tY/+7c2Ho484aqOJbA23gs9+cmz4eGtTSKxcrqRYiHo5KupLo6+my8zr
byu5LNpa0wqUsQRagAPk58zjAJYGah56gW7W5vrHJo7EjZZOUXquDRNhcCze6egzYu0o1cP94OyV
wZIjmskX+qy8+lUfNJn5G/skuTRQ6hCBwTPoEFsZnHXUji+bKncOCwT99Su2t4mRw+oEz04QoQVK
U4t93oywiB3CcXOjWn+qi5K4RQ4biYKYfjVX1nzYMwWTiLA0Edwwdfkn0TiWXMqDqUt1DiI7fkxc
uoDms7wNeFDx4TgJHIi8HootmOdWvCvofZtUQnjoCXFXbZtVNthfqhiCUmBy4/8DPpO9abgh91Vr
I0UZFj1jPWmS+JHBbgd2y9fpcUQv+UI4iYz0ok/XPQZWrN9ujB7ZmlYho8sn2NHJX/Rj0i2EaxqJ
beEKAkwyKHM+i7TSMOnwAtZovr+kAUBoADo+h27WC/GSeTtpAgetDXTzwQz5Zlme4bBUudW66al5
q3MzTnZK/ugIFi3e98bMJY6vyYVlyvVDJZVK9EOnhdNLA1UZBG0+usd3e7H/EPsm4bt5s4/fo8Fn
8zdS4lsQ6zXJTGFrBCivPsJyXj1oS2dggn9IFq5UmdSodNP0A/L0auCAlmHYKWFwoQoI+JZPigm6
eFlmRqj8rbjY1QNwqP7l8XbdjejdhVMdDC4J5NTEvhPEdiPtzmeLX1O/sB7azNXM3cExfZ9BJoFN
72JmaX8sPFPNKzlyKAfoaiuFQfT2i4gp6vTU0OiBB4ERr46mFLit/9MByqqs8urBuEobgauYL2mS
afbb3uSK4vuytdcIdsWx5GYdJ+hCgPpGj6feHLE4p9AkzPuZoS5yohu4KDmIj4TaoEMHLmVgbuMS
F9PrVblPZ19T4GWTj0sf3drZvTMfxSoAtT28qlLDfOAQHKF+LLNl2d77aZJ1SeT26GI+TM6GbDn0
JJFZNPGOsd9YXj6q33zCvGDe598KNI9/LJI5RnBlyZWdkBfPvLsJnjOpHU0zoUhv4EkI288IjMy6
3UljKb2njj5cFXiAj8VyhXl7U+BDa5Dg2WE7r87MH3EePTI5dwZdcbzRrQgOc9/N9C63kT3fP2wF
vRu4CjC9RCMkRh2I2b8OmhU5/eReM+hbMBsyiyz0WEzCWz5UQXo2AM/L79xO/wSTMHuKp4N0hKiE
uj/9LabhTWdIrXFirpnVtoebNU0GNBT46RKC/dJn+r9hYQ4E2jLV43W1iXfhO7cVlA5Td4GI9iSS
fxMy7fFiheGMMYvKILT4xxkebm0uetq0N62Bk908lmcnDwexroYmnnEmvSX6imGIluF3H205lW6I
/yCuKXTOr2YuJSJpzsQZnQMH2Rkca30VymWpBWVpkw7O8rwNNxUECmkxyzKp0lwaN+F4ZC0x8vqo
z/EMxdtLtDC0RET2hnUxxzvIwtCBCR7+q1Qnnd0lIP8w8jzERWiwGXlGHyHe6RJgyn/g5UgBZe1u
5tKPFExrddfOeu+vp6Z8OczojyYGu/ywr5AtOnWLGAa4gP8FDeBoTWT7ZsbOTAo9hxGrKCo6wfwg
uTQmsoarWUh5KVjEGlHR7eTNdcYj4Pc90t+SnSiW5STK5M0fNBf4kvr5OKLCkEHF5irfQMjH/It8
qFSH+HaENCIJ4OVJx4Y/FqABJzCE2mBp48ScEISo1woBLjtZJS+6jf+xcEeMwlJ5q+Fh1RtLs7Y0
F72zPsYVtt+gMXavMzNualo8nq3IsfYOXoaj8JrR/XhGULVng559lms/evCeosU+Z1v5SXVLGxb0
bF/01kWWadQYgrQrwt8YUHCwFuWmMkHGmPkr9di4lWtOfp7bgHaLeuDS7V+Xa+HbU3eIQYzV96bd
VMDVFqm8SYGIE+4LoolSoejH3AXdMjCnWL9ACWUNT0hBudp8wng/b1pXkxg+EMElVsBzRFc0mIcm
1neDLrMBjj2mhqL6aOYjPavj6QK926VnzUppM63svP7Wvpt/7eA5SjChsj4FInraWdUaeFoZHss6
bCjGio8a9sJudpHfj3VqzQzc6yRRCtq6hh3ks4PCwuxwC8RaKqvhvVb8a2PnBJmEb0hTA8Jhw0He
s9H9M6oK4wL7lTbWv/qrAXSCQR0j4vhNWBJ08euZh2vIKfcmeTegtJl4/rBhwDpOobPLsl4C0XVN
A0g4pCmqwsaR/cQJu6QRy8k2WMnhG5XY10tnkfly2d/v4o0Ri2ESagGVjDT4bFtC6ypof0UkLwwp
VJOA5sFihmsCjJtA5//tOpfOWp0jxUhPhJaIw/Xs+Ba8hTrt87/GJAElMRAyliTTS8S3+gU6zgTP
oPTzmJYuPwcQl74HKqs/f+QnaXfvFhWg/A2eSHX4vc0pxQc7eE2an/EvMuQ2UgPnkRIG4NhlKOUn
uuXMss1/n1zclXUkziYGYApvUz/+W7M+AV8tQa1GLz3XK0vZkA5UgzzpaJPSyxdNf39KhNR3CYIv
Ky5vhgJ7ZrrwtOJmNGje6qEagAoIakJAP0C/ol/QzeVBvlyWmghS9H4BTl9aAVHLHtKmtqh/Z56v
BmWIIJQgAToc85M5ycWZU2DjaZtnVTVZ9KfFUkHLhq9XkfbSezrg9670r+OOzMFyWo20lhBet8kz
sea6zjw1A6ogOVruP3utynWrOTGYT9tpup/qYbk/R0FbqbvnHgtLOFi+3W646OOfgjAqIuXaIDR0
SOlqnp+OFgJvugB8vbHuFiOpVil+dWe7qIBVC6KSY4BM20il7vQifNElATrGO7W2agZT0UgvukcB
8woQw3GOIoSqCoJnIbdR2YlUGuwuJUBKmb4nEbwSaiVtx7/dhgjT1dLbsSeE48+rg8d1vpDMjxQY
2kdnHbrBMBt6a/Tx7rATNkgKbFZ0VAXGX4N20Z6/ESbg5qIcZ428xuuVTTjskvalAv30sBc0cqB/
j1R3ceb+JspDH6xh6Z4CgGq/fRii9ZG83mNhzT3++/1tTVjk5VJb0XQgHQBZ29sxrMEeapt6j/Kd
6sdKtqYeREZRVgVQwtv6gawtPanruA7B89VZx1mTS0OrMeOl0zoD818ewemop6o4M8E9raaGlxWB
eKxZ0edJKbLkh0HciSdMN/1lQY/YSqZjjMOsgoZZ4VFnV7BntlQTrRCXC7XPWXBJbeB9ROtB3ZnT
MsedBrQQ3TjaBn5/qHh/in1Z2DT5fymkqs1aNkA6cDjELK2uvTtTm98RD3YT6en/3PU/e04hkHiY
aLoE2Ivcpry8FTAqZkXFkYdTAguu3eR4oi6xN93IapxsEw7QWhD9WOGcWX9tehXbJ2zIJeUYfAp/
vChHWhHvHEiQ/kSsosj7LY/rulPiI24B2/GNM5jBLiyhbHoMkT6UgJHr44kN54vIQfbTXBHTcjIE
nuKdmwee8scfvcxZPY9d16IvcafyvRbuDQZD7eZYmrRuyowrUHXLR2ZJpDGPEnKiksXCnKsq8R8Y
i7YS5AwREBdysBcb6eT6vQ7EY/w/PawXDSQ1m3HrQMgLp9aFrDT8P065KKT0cq3v2oMz6eGQOw1A
CrFa862uYXCXPMehZkvYx5E8HbEvompmrpkfQv1OA0yLa6XkRQjh+4G3s3aYpujX5EFJMls0VIrY
8rFKyl6+H+kwPfUj1XDrZxbwtKmSA4E+z0OQ1sARORFe4++taD2m+HS3Xign370TevAHhkF55asb
ixcBtjNtsUlzj+27ATsRc235EHfEhXMBEHUsNpNHYcVappIU853w7Dk+OFOIaixCTHcVV4niK8+v
fxsI7R8RC5vk2RDqPpUFFBZvMsSF4o0HwWsbrMwqFBvssn7tXSYcryRxwc7rvKEzTl8aFj1at/hd
joP3wYC5wF9phMiQ2RTqzhUhJuqX+2hcUBu8rRkJzmg0trE+76GMHIS36YIVtYLEBtwTOWpMEq1F
WV66fEnzk2bj6X2Ov8DlDLTSqKL5ZBQ4JgwU18cw8M1Nu4lyXzGOxC5aHb92X1gb/6oUUXbi47/r
i9dzH5WbVAUuT5lQFHPZW3wbjvjQqAtZYwtTmprYosxPHUZBrDSumnhix+ST2XZTbFBuw1kD7QXr
cuopO3fLt5FdzrRwRQhNKzE83FEiCN+xwVxe0q6dvaD+AyjOWEkwE+KBIcC4LiVzDskQ5CP1uNHz
V+VDwWHJ0vNa1WrKVwunelDeCIECfWuVnbz85lX7Lz83xJkRyYwigie5KxB3QLCpvBWaIBzVcZ+0
mr8qfbD6vP8AThBIuleRCIFmqIr2trt2EW7HVbu5eKvGOPlehXqJkLNWj83LV0BOq1VkqaY5rezm
g4FsFYu761dEl3bQ1fgz3/4wJ6uTS2/qXqqAClHC1rrhxPFZnz++iLrxsHzx4GDmT60jZpVKUaii
O7/SVzy/cfqYCuVa4jdgL7TcCZ1pnLJGlFxOKTxt2iSyfGcup4v7E0eYfHhMjx3Be15C/IaO2b+u
2XZjZO3OZJBPL0LjQEJMuqxGzlTvLjR43Q1dQLDeNE9AeSUQTXEPEHH78+dHgeaJXpZG7jdBntRJ
g/kKlVwqyIiLkBOttuSsK58MInnUy2aeqyobt1ufOym2abr3/E1baHLn/jDc9+Xa7/DztUYbzDEB
JF7ZvowlZFFdNMoxTFF2RoMH5U2H3J2tkxrC0kNi6Bxnec155OjACxPO70LfLyF5I+JwgWegWZmz
mxSUBZFU3DGa8c0uUHDO/A3EyHAWrhJcEeURAL4JJQ9xr1vphlMYmBBXO3+HRabAenMw1ptfOoH7
l18adlFpk5YjvhNvLmpXHUsnWLjkGuU0WiPk2vn35gmuuu/1p1+SFHbxaMD4aMAouEX+oxvGv6oq
UJlwytnrs2bKKe5MqZO4Wrmb6CZgtFZvyI+QBT4KDjp3OEEpSNlBuSouaU/6KoVucRJNU6dSIKa+
swmOgqYloAakFNNl6l7Ap1VZDO6B4E7tKgeTiH+SUPkY1TjVzMLm9o6tkezrA6UPCJauM4txXaJx
Uh7k9LGvNaA7cBdg/HLUzTd7814f1plhR7gajvXKqL8PbKGntogWCbfurjWvFHythLe878YbGct/
DxVrYN9vxbjOQ6pEpjFUr3dRSHnY+Q6DD0l2tpUPosfecaRCJ+u0MdSMCTAi/PsiiAYTlxv6yin8
gaIApv4zoEhUMx3n/7aj54JO95j0ZFa0SLE5EiURXFh9mETBWCP2f/vNCNjBcYgInKklXjb9IaG3
Hh4z/9tlPoBSNQM1Z2QjDYWZqeaW/Wdj3Mo5xWpE4biMyp9jD3kpwGx3P/u42sWcvcFT6WXh8r4P
Oouz9HUoh0TMe9IvhapJSxrEOKUQWf+9NDHSvozomSa6zNlpx2OJtzWKPMcJra4zTF4xsriPIbWk
gl1tHEHI4sATEH4UOpgXbVXEn6uWlw0pYJxNsHzmbbsiBSUMUwRB9cBDlu6DMEF4WMkL8Mcz9t8u
1YIAvwfdi/fpdrGADpT9tI/COEF5qfiABXFftLBvXU7PYDGWNVvfNpq76ZrB+Gvw2J2f1jMgxvHl
J5FbW9qBIE7MY7NYULmUmlfRHeytE4lNikaFDHQrxnCCg2LswnU2NRtENiru30944IKUjlQepNys
7X3jWPNVluBgVOk0hK1nt5rIy5iitdTbbMTcvgO4yUrcg/SfkQKVZEFPF4DaFeWR88El8eLeRgm2
z8yseb7kgPhMt9LiWJeEG4oGqopcfFjpxVH3gwEIkAd42d3C4wiCuYbxw6bhl+y+oOJRXpa64G9b
LfZrknoBlLeoGEHCtUoK2bi8iKeLwq053Una7QP4cx7KUCQinNw6Ur1Bu+LOIPwZ4OhKCZsL45ri
HByjaNXFbJ843UX8u6dKRE96SO+8nAkAEiGZixxqBgWECLWxVk3I7j2ewz0qc6sKA0SjwQDP95h+
dLlIfnekRrk1q/JlXnRwnktDzvrOvUvkIN+E5E42QPH8jff2zROboeADGGXy81tB6x9YZqVd7VS4
hcBY9OFGOQ8STHRSQl6jlA2356wWf3Yg1L657MaLP5XdFa67IsBibsLWlzSLgPuFdqE5lyPw6Xet
75tvzkq+F6gbv0BLpD3lbNwdkRSRxZsnjUTOpYTlc2THMvjPfIbdD8gAJmM2/DJ62VKBaQkf4U19
/NeHz2mac0yhL3ESuIGLW1xzXFDuuxFpnqnMR9RiJ3Kpc+adiyQ12p0O/pAdenzSkyi5Nodjl8/Z
eb+NHVxYtFnk6Se+3wjIwP14oLGsNnLXY3cUEujFMMmJMO9aL2+VInc7DUTnPkobjmZxrUsGKf0G
DV3+LV/7FA/8gpiA4p+EhALAeMSDubaTkGhFCF/VZMJvKEyR0ghxztUVHWLNNeigpc64suuMfoVi
bmfvZqzu3PYJSF8DR8akN1kYJIgc0Si4y09Z9ZUktvnSI5+tSZEDMP3um+O0T0G4qqaDyvqwiz4g
nDJyiIA9IYB1Vwz92iPSthxGlPko4UutaQXMc6/Ku7jfR1avstVl3Ay5VCfAfYa/pqoIbg9lKNpD
B+phZjWWoutntJ8ypGvDwQSRoe2fcoaqeq7B/v0eo4CaUL8Fw6KAbafs+bqRsV3atJDp3gVLIbiU
vTvlenM3i7zcDfmpn5Ec33FqmNTTjlqulia7j9Zwo9FxpqCQRK6PiBLVIjpjM4XH3SNo+Ml99Bdt
vEwTotHLKeraKEqRcQ/PLSDY4z3QNXYKlTKMF8yDvVauEJH1axErf4OczcS22QRUQSpRpPGIxB10
yGtGM4ZShCJDXyuDE1JQLqJ2FyajajCLcgcTRmtxRQD/EzlSyjSn3gAFwMPSGh9DB/sY+cgYYp+N
YGxviV+/nC5efeEtvABjWo7IrtCJvB2QSi51YtD/ysbY4/5ChTuBnrw1U06Kw603XWaJaaEzKZn6
YvqGG4vovFqWhQBPKn+GxQwjDGCDO1n5xHWpDdqvEAWqOf2cqwmqZQgFlW0DGtwAguJG3aQmtLMG
wc5rwRwn053tUR63N+RqQN+mV7rkqBt+Cd91z6ejbr0VhqXU0SNMs3G6XUzg6rL5gJfWIduaCRmt
kA6Is6wwuM+iTjjmZfhHJtYkoyDMjcwoGGfnr6gOJ3VMLa70A3r3arDMIKeAJKMqb5HmvGzloG79
7ifxFfXg1PUuFiXmrA2IMM1r49ia6CCpY65dLgk3zLCnXXuGdSOAtC9TFS8fy7PM8vbebf0wwRuh
Q+/jB+thuXIaHgMkgaj/EFRcqg5kdKBU+bcfK1PJ4yloivIBPKj0uO38BbQIaaAN3B0Kxk4GDAOL
WVOka+pZ5UkSyZKhhKHd+3UQInzMOnNcfZGmaFhjIrKCNscRs06PMBAqDhUS0gosQAQLc2W5AQkl
lEwJ4xBQCz5vooKvT9VP1ljDzvBecbUBnt/tNgcdAoWeEOS6o4JgTN4yY3/GETJPhw3m9Y78/pKh
mocP+mDXo3oREN5+JA3vAEuRERPjloPFF7iHYOaGc29rh9rI1oJvWADJTU4+F7dRUGsQ9nFtaPhF
dvsDL1RkX1q/cn0CKydWGQwx3CGK95dWxBv7ZuWO4BPMvKWFKABXcPgIhCJAytTDl3P2Mfhu2wG/
XFWhimnuFezcFlylfjk8I+7ZTgIQ3zxKyJiAn36LxGwJC6s/j80z+wFjgU3NQVaB24ON1ez81SbQ
j2EwfxV6B5nhTRldWoowRQR3I0Yg7AIAwqqtgfCHxmKq6eV31+zienLcrKwi2Y/9voY++G1B91PR
DMNCNRXqwsgFjKZgOhgstq4R5/2wVPs115+zhTSwR82tI5vI2LQsHUfT7M/2WrkyrUF1NqOw6oOX
fT9eeB4C6/E3ApOojBNZTwTHeU4C2jJpLZ8LaLtKgOozyJRZ/EZwQ3H5S1kJs2Xgi15Bu+YLKLGw
vi3h5befZeOFSY1Kp22ZDgSU6XqFhaAl+oYiwWqH6VLFjuQRs0xzugTm/yjb4l8+gAd0gh2scUYH
qo0iQtxF/1z28M1uU2z/3m7DP7Y6c0QJ7bKmg+kLirf3qhKuXiLGPJ1n2j+CDB/x48pw2xhs3TeL
AKZAgSnpmEJik9ACnBCFevUmIrOAuG5CqQxOHvx1IRt7jUZnRPIc8nNB88jiOkW0wmu/C7CSdjGu
Z8QnS6GbjtNhtk7o8yF9GDzadTlaUPnOKwdinUbcc/0A2FGZb67LMQPkN4MO2BFw6aksn8/lTzo0
IQ2M9nmF8kxYb7j1QRwpXjluw+3B2ygijZiHE3iPB/QUcDkD2IneneOiTGyhHovI/H0bsVRAjNFb
aC336aQFB+BSXG3ov0ln0t8LdXG0if/tnTSFDyXKGBXDlE/yUaC6cgLkYPnDh47IGX8J2fYjBlYF
yiZp1DLR56sIZArYJn+3c5avpAshrQfenHeRXjYBSCzpzRf+K81dbJ7YFL5RlqMFg+qEq0e81WuO
mX92nIrG05yyehwDDP/lJPP/574M0RmWw3c78N/nOvgZWpS6PP9B4alZ+VC4fyUkkblX7S1ctNcb
gq46utA5Z8tMSGZL/CrKqfeCbfL5bUUHCq8yni4tODYDomoGXN/yInFQYjgq7gF6Wg7C3MUI+Ct7
/OnlmqaYODM6iK3eONy6GKXvYiaVojP3D2zkY2ulRjp8DieDFl7hAhweIyFKW4iLk/NspGKNv4QD
gKrQT7RKoc4ZmOzslTuW5h6oAASV86tnIIqwq3FO1+X1pOzt0aovJ+flYY83A4d/wovglmSalPg1
60YvyORPtzlRzR4ayelbY9jwi+hsdbJDGUG9dKt70N+I68K7gDsHQ4bsMAL9s8HyvUX56eC5EHc6
tSCxjwT8tNYSzPE3h4ZkX3w2yyP3zx/JQJ1tChzkt/ui8o745R7SivZRe/mhx/c2FFo0LOCgPtwO
llFv0U8whNKgliE5LDIsipcz5djnvNssTUJKhJwQKXdsNLk6ISt9I+FmOCoVYBg3cw7RuGQdzls+
DdP+/4I5FQINh/L2EPVYAJ5ga1CsB+01JgBys4jjyNHpYkPwG81aNOREMMAPYHqGNmFo8XwnMlRn
M93nmfvWmbAVhn3YSOOcUEMecSVG6g/r2QSH7x5cuae2s5HfwaRJozAXOeM2tjimzim5l1Qas/LQ
C6U5rWC6T8F0hdXVmdZeTsq1mZA2PytsPX16EG+A4EJWdSL2CxkC/W5BnLgU8n9mRFR7gA+C1Lc1
81FTqZ7TrY0VYOHfVnzb7/b2bs3fhOkTyFj4IEWWAOvlTGQTzvkZiblmmagYD6fRI0mcIGpIWAy2
AavDc+hsDt/4YBS7AocCoL+nv7TQEBFsZjhMbX3QEtXv95Myyu5ojwKSl6o9+wjAd+17e35eAXTf
2yWNN/KrXnvSdG9VwXH0kUMBjNVoErxixzeNLUr+ol7w0ZL3VKUQWfBiTBcKdNTWaRv8qVaU7QY8
jB8J4riNCu02lHI5eZjeN5WTMu0Bk56YMG3C0xCGtZj4VGNfcyHQHVTOzLhKwz0EimSyn//QrxvO
WxJy0grabOwCL6nYCEYYEF1lXREJMa7FnhEh/SeDij/tYnpGHieIPkHhQ2iUR9huQdcfj742baX3
C8zQZziae+uIJL+7xYKMytW4t/Ecrodj9/v9K5Cko1SqTckF4N167IapwSuSkxNz9/JnIxWuqPOK
W32gHxyw5gmEO38/+QKxU0SV5o/YAz4iWYQAIGnNKVGqyQ1Sdwf+HkrIv2lzjYO8a73M4bku5KK5
cIvotovThBv59O9xe7iT9Cn63dZoaPJzmkjVds8rmVMCew5S3rr43ig6ksCYVZTfRdxM6aNDddJe
68J1Fbq/Ka4haLtVDhJ6ED1lVm6pmmx9EIKwyjv8Fzq/ClSr5QIWgu7mM5/wJAxGz7QD8w+0Dt/o
AhMS4DulpBySIC+0usR7MRuJv5ihkcpT62BCr0o+8PL9K7WYTtEBVxWshizOUiC3muHENva3BBnt
dPFgwgw3/jHUKKCeKMVb3pGgxuMDPAUAgiqrOyvFfymG/S1k4G51er/5y1BzwAPc/qCrPybmUP3R
WYeEiUu/fyQS4WUxigk9J1nzWcmDl9I8dA13tHwtnVYDwLlh+fThxY7RhEi/TJUYKBo354cGUBub
LKi+LrxiDAcFsIflvFNS+cRXWLnLooQsrPoV9/5cEYRXjp774t9QHiLhoKtaBDQSYrqyM2uyczao
XzVXXdWAfEqLcXdi8jOTNQw+DHwDIlxtHfK0lKQrV5/qlC1HdQiIOuzDFNOxdtho+Gh3dRSUBYIz
4qVzhExmK9K86WKD1TMD4wxJWHEYCHP3/tby0DwqTVcOjlJ3v02PYho6/R2hhncwZU2BYdizbg/B
rwoo3awxHC/rs/vluqeQC39bJU5KFFk7+4qcHTKLYWP+8P8iZMqHo36+CCrITtr9n0eT5DvaMuJ7
QTZoEqxgaSa21e/z8XrCVukU/moF8fhZSHWThLvE67bcYC5xHnJAc6bPHILKGMQN9jwz/1pBEkQN
jM26nI0C9BM6jYpb+7WygVQkj3/7oaVSwcJahQ7UjjB9+WrDoZbDF717cnRfqKXPrQJfIzsf/rir
6cDO98kRsR8UTJ9mVrt5evBVfPs1U0Mvaoo4fA4M5lNq47AkItr2VUeDVcrnlN1drfboqIN4Z19D
58HqrYGcZE+B4bhT8v9qYpVjLd1IP3HcCMxzeTrrRg4C1L/8JMn+keQ5gGIfeB2W8rwy23YuFRXj
D8YJuefS9P0oJojbP4ibiF8q86uDhGaEI8aV/c9ZBlvIpdlhnfBvgM9q8D3nJhUXhFyGcfQ3a1vb
qGDlYt5ezoVio1Xb27Ka8Q0xTCdXeY/kUZW/UIsg92lD+Nw4ZK41SVd9fKnWV/6j1l5Xn+sz8fWt
l6XSXf+auWR0BNyrmNCrDOTGSKjEz5gubbynG4lOUa5QON1okFg70Rz+QrH26twX7KHf8Nxe9+yU
D4xYHKP7L3tW3+5/XMOJbAFBXV6Cl356HssvL0QOWxeCxGG8fD1RMQ4F7A2xFY2YllZhT9c9aEdJ
mvUrZEsfuyvTNLW/5LFzQOOlnLWSu3/04A9dxWQgwUvxqrC9AuWxR5m16y3R1Nd8kqZPN60vCqtg
qaN6QPoX9+u0awg9EqHBAlhuwuUUQ1AEkxDcyuNEHRSRwbMBdk0rhkR/R3MIlME/ny/2NriO7Twh
o5lVKTUmJ96nRKwxqVJqCx0Us4/nuXmR1JQ+81Zjh2eSYqWERrSOt5BPJqz28ldDHz2SxmLyfLoE
PKChOP35Lh9qagXaQNdgI1JiyL33CQJtlq9Wd1EYC7EbaehlE62Q7O0FhGXO6ugdE+KJUSZ3H+o3
q0pRPqpz5Poc4uEROQWxed8gNiVxUhpQN4yU0JPD3I7hCCH2jB+vyzYXYnWWVa1LiXHB2zI/iIaH
OfgTYk94dW7q7JbwXd0zzvs/xUYxki/J+/q+6ZGgcfdBQzPtiF9YXbDunvcLadOWVkaVGAgcQapT
AOGISYpi1xXytsueY9vHycAXFPZDkT0NmyTb3sbXcO8en4UDDlTsucgE4JX8aRzO/QRbV8Wanks3
RqSf/Wavdd/AtCQGlxa5VGeVeuvBDZKL1ODn39tZdzBPzDCmt/juPe1Bq1CKrt2sgXAnBFkzwI2w
uRLRGronTQG5HKzhbTY9syGebq1eRhijCtqQfyEaSiaLM0FOHCkXwCyETyu+9GeF+69g50jWcZKm
Hykeb+xBAr2B5xTjmlbhZdpfyi7cAsRmlqzVmA1pR8y2FO3kBM5yneFqBN7Hzwoncv+6tT0lnzvw
PpHab5/iJSFd7ilI2cH++qaPKJHUsae9qQT2NrwuS5yMxmDZcUJA9jWMJrrW9Qhobw30dAv9bEkx
qDunPKbXnlhs7Mg1KVObaLWf3E/vxZRtuk5kuJQxvLndJm1d+rU2a4IZHTZw3lpFyNNDIUJ2R1Gf
RsZKLtxSGuRHIE8qDk8OUg+niwYz0lq4fKEsDHj6VqEhhlL+MVSUOsG+yInQVMD7rIEjQqpk8jpn
FUGQYKoUiBaDcKnng5aBLZvZ88GRzn+yLOeJIh7x3agnqxvAY8ikdY8kJ6MAmItbsq82NjcRdWDq
tMF8CHBQn1JJN98N48x15Fcmd9Kgxb68i81MU68FF3PxsdDjbF/eWPfDZWoTyEttwHglEAUunjjK
E0ckw9Ps42aXaNf7yTn2EG8HTfc9UWydlzcBtKnLYmUgTKjs/mzRhvQSP+IWM92EnW6JYMZPahjp
Rxo/pF2Ct0cxcR/uowb3zzI2FR3XtSPkVpr7O+7n2qaZ+Ot8KxhYprWEDT56l2AEs4OaCjTT9jmB
UILZk76X7Uigw2LL0nZupFY2aKzv8nFthe43n8qT/rW5nj2s7u45qXokbUhpi4VSUa1lA66J8Uvr
G9B+yhOVfGf94wHyJHWB3ij0QUFXh6xKITuuEi2R+58kGydqyCHK1AXK3pKSRfxMWCy+bdzZl+Ro
6V8wwgJdCl4pwyRIJZ2gTF0jji9mveQ5wo2oIhnCGxiKtwls/jI8t1RyhtWZE8GYIBwxCQlEN84s
hvrznos66GsNSCcx6YzYrftZKtFphzHOPLY+q5b7tL2994fL5c7XSGN0NVHfxGctCApE2Ebf+VTJ
qvm9UI0BMxoJ3O8YrHDO6yN7ankVsPBCjh5UiJr8JZhYEilmw0WifPoQTqEpXX9d8zvJkKRMIrMi
sgrykYFm3sJhLubXibXuZu+cgd0DjR2t7ourKJ9rdUW1KKzE3U+5CiY2n+enGg+nPa1kw2QKeV2X
4OiH/obYYgMs5i7cz/vNyO7pVuiXbXi21Xrnf/IroL3bNRBnqLqjVvWAlP1iaMIfVGsg37HoWF2/
V/IH4qJelOzxb03tANBp5izT2AQT92lg2oEtvL60So0uifXLf+gXBo/gPBygoj0O7swouq9Rro6T
Psrz/4KmswRULl8Em9B2CssngdrOx6Dnq7+GP03p7B7gotW2qdiXPMT1oWDTsifLCXLSOgDie2U9
3YWAF95o8IduxppYf7pn7RAvHwmN/eDKeg2Cja+rv2Zs91pQPKvLIALnlwofe/YZ6z/5FQclmz+D
gmM/ze63TJdKk2huV9/N4/lrURwqjbkSSz4ghcPcpjQO+dJ9tNo9UbYjWlHKsjf/RDgCL8eAm8n0
xWGkcVoLrJnv0KIaHTqQKDsc2rLwtc8rONQ+k+b1qUzHvMZDvm3xJHT5dId95v3VjqsfpTfXoqtc
R0TibEc5wk0l8PpkvVHM7nLFE1SfiVdwjmueQzqSUlTs//RlwbDdNMsbPz3DbZ7p1y0DzQ7rE0oD
SQqPcCvUK70xYjDZjDkYRJlnctm9OHO1cANdnTAoN9Zu82G7mQo4GBL54rGA3AV3tWPhTQBXq+gP
u3hNknd5R8+IwPC9MhLNdaa1wKBlUrOOkYvTkdToNirhHR4MQYOSP0F25xxLcxqWVazGj76Qp+YV
HFeoIl/I0kGUG8cnMYjY09N9pZhKERYBH/agsX6IPJ8/eyyDPZkBMEo4jD4XKS1/gu3zOOp+y+J4
Rsx/ScOMyub47URCbTwXPhDCVECBy5wLKp1SP/W999fyoYntqCLC4nghOpBuhKU+cy7LAgMJu/VM
Hn/DAoIyhdogU41CFc16r6p77zIQFjrXN3QUZ57Z5qvdUsmLkqhbC5IU/CL10Pj5aUPupcIDikX1
EQsMfzM9FBud3BeJZ6qwOWPJ2IieBjnjyvNtn2/4ogVhsyZTR7f//mC1Er94gvg0xWlMj+XFwacE
AfL6l2eQbOH5E1XPqzUwM3e7VQGjwgfKNLZSW8sjynGJxM2WGVGZpAMkiQ5xpvilLZvdr4SKRtlJ
jjgR5M9wgIQ8NLMUbzyjcvmXfG77JpRADdPx8EF7qHzP/JMEQixCpqgKyyR0dSJbL7AJPMEqlCyL
4KjdlOnP2gn8qZ2VcaZkJ+Z612F9nsXOte9EgcBJGjDFs4fKLoGtdKz0MiLyG0h+f6wPO6RBdzPC
6ZiTonHPyfs+wzn5HQfprfFSmJLRzyTQxRfuxJW8UKZos+fGauC/D19CSiRjsSrpUMSSgNgXGNkN
Vj0eM/gpTB39SIDdmAwZEkVb1263s7wbbE107+2+54z908oZtRGpyaDrWZ1wJu19L5KPPkjzdGJB
odFJd7DBA+h/he3MCJdLL/bOno+gYASiYbvoFoGXVSSICfhlRXGkhKHvaCs49oVJ51Y3MhQ/GhR4
6K6jcoJX069v5pUaupLGxfHye69yzROcQsIVIH4w/kjKakJiCPI157u3hkwokniWlWjyrNa+Np33
Q/lTtO4j8v9aBWXbpBOkrD2Z878IWhRlqLQmOKTOLp4T8of5toD/EuYFwUMRr7V53xlwXtF1JzZ8
hsHcwzqZrjaIy1jRk9j2bIWqqZFrj4kAto53F4vZpTO+jX6O3fY23iDtqHW6Dpr6g7rJXdEiQxRa
nEQVP2+Rob2gSHT/lCVdmU9V/91oh3AW7EQjH/m5CJnqOGwPSqjCKh+oHWp5fETXaENo9chaMRya
qOv9FMU1ZfetiEf1Q9bcOnGOZfAsZHV1aBqDPQKF3RMdoJpajZBkrR7X6hIKJ7bDnvMx1ON/mpfG
LzN/gH1EEmzk3Jb7BcSplPhv2qHTB5waVhMIh1rhC+h2Iw7ZExJcjpMQmmIlouPRPcHy/2ruXRt9
HPcwqx17uZS6wQ/SnAqnTmeDbYG8eyFT7OfsdimcBnZNV50Q98GmfRXZQiDbCNmD0k92jX3epKq/
dj2ULPGNHQSDP4S5LvDF6ScUWLyoAGU3gK/N0OHJ3E1q1nyZ/wEeeSRkHpiOB0nldWiC438Yd80z
JqMxY6Ai82RD6P1jXu8sfVfrtH0BIJ5TSQW497GgeGEM9tW2DjhZRote5o0aIyO6YsUfoHL7ZENT
j5g3rZ2masSaClsHQ+3+bSFXj9ZWzmK41vLLIVYeXEFS73ypgkP3KxaSVh4NbolDTZ9VGhkgKY8f
baJ8ivrTQSNmsbkN2sdcXfxMR7WVOJGASrTKyi/Igquakn7ZMKPiVK1rrfCBYFyhIN9amxelJ1uB
YRHOnbFdLqXIKJQG5wTVcpllJoT5LuYJu5NK3k0PLHLTQteVisT5pgN7OVPX1Pz+igmAEJ6BRas2
PPDiW/82UlLOCvm5JyrUsNa2bvhPxrkXdesg3VIRN3/iOxwtK8X0cfu0ou1Vo0Sw2JbjHEqO6t2N
HRyV2aX7YSKqPmjMC8YPtuqjyK+Mzgbap6D0ItTigDpjyaG4lceS9N8YD+E2N/gmG6XrzBI7DMEL
RbE1mTtPZgJsuZvhVewpmeVqa1iHHuwhLkysnEjtowLuQ3wJ1Qy06hoypKw/cW5aOZhwxx41J03x
hWMXzDHaIhDH9GhnrNi/bwmrj+iyTvWRMBybCwXopaHCa6SNjULYTBAEZbYdcxkBt6z5Xiag/Lye
/mXVlfK3vgtm4o7ayByuTI9JPFxSp9uDuYu5+ohyZrk6AEvIcC2t6Burol4QOiwSbosDbNyq6iga
dk5pvmlhtaG+yzDrH41Ydf03rLnGJbNNEpHKx4cqxbfGyqGKSu4RkCCEpTTOgyAqEoAsdt9ATQp/
GjKhlPC0NeZ0QIXnRMuy7pAJ/LcRGTxoMFSvUkjw74N+fHmur868+Cajf5TzPuOvUzetwHjgp+WH
g55o7F2vCtMpC/CfYvgiCN8cixyqA/ZIp1RzJc+gLZ+HU1MWcsuc4AulcDdhRrkOVGhCXmoVTyeK
FMTJBRL7cXaqBZxGNoSn4a5d8mEacN5UgM5JtppTTVGqAx5lATfNYSXYv8Os23+9QIIAK9Z6xMlV
j/7Tcx62HuAe0tms6EZzOpGohV9Myw07zmPLUnjRsooCjstw4kfnVYq/cPRb9gmj7ROeucbeNKIc
YT0egQckFV75k/bLC6MhjTBkUbponjXkxtXsiI0x+FLH94XdeXrKVqqmzBnTtSmiSOGdI6dI8tyC
+H68ExvavaIPYg+b52yhRZlENfOTceJjTzm7ksIXsoYybzllnUNaQAcQ8piooVskGVJNS0u4tRGi
BBP0EMbtkSoZn1coXyJYKdEF3rj+dxJShan+ReqYAfEGFE2IV4TelE+ULjF8HpUTjVspnfDFyaiv
gU7f47ETLE2wkAnVTLOQrSBAhwSzRJS9kDGgDan9Pi72Ceni+D7QfUTvy4DU2I1TBVnjfr5kEpQb
bxD3hFreFqns1VBXhzUWBvWdtQWLYQtV0aARV3ah3d5UNko7KPbX7IE/yfwNgRn2MjHuCQ6e6HUr
6qatti0L7ervG/hRgiLqjn7ox8+rWLga2Ajgqg28pwH3yzPko1WVXVbLK53wC7QQYQEM1DBlGmjC
q+e8o0KaYIqC4x8yuCwKuuZ81RIDJjYtk87A7F3cDtDMfMAZ0xP/gRq8X+l478KV2MAavOK52j23
j+pH5azosGRyo/mDpudKWXP/je7cYOXoUDn1xXY72aPjWgAuzT+yVlchrfacwA7veU2+95Ud0r+D
qibavqvuIzve2Q/cMTS1gFQxcsUnxy0VCn315VqqkuyZk1+soDJYVKxqYE9UCkt/+wFsfqPHJzeE
EuEvrUfpGU4bHOAroDhUiuzgqBTN/MlEmO0zDsDPuU4ZsamKR4fDXYjUGwzW+JP7Mkuf3wQIkP0z
cnvxt1ZfPbvnkb5Eg6pdL6x9ujlcv3daYBnr/ntQcQ6BIvyXSwVm8yN/efhC72w15ZxcKJnjcF7U
DxXzO/tu/Kd3cD+aB0g6PWNHyRTx30kTFAJK4oLNHkOob3akRDn/5CXPpki5VdZzrZOC8HAT8Xpd
4oZUivRPUk0EV4SGSz0PqPq5sMwWj2MYRi2diGGifXPH7rBj2Eec7/38RPT2RGzo/KyqSMseTIjf
PCT7FW+NhqnYuQl6t5zl8ND2r2EXBq7AMVTIgEZlNWl915fqDMJWeFlShwlEQtiFB4o/0fieGkID
DqHZ8Gstlt6mNmz//JqH7Ub6seJPjhTRGQtzmVAvZpIR9HdGg7jnWpNkyWQ+xZjVUBLY5EikySi4
xfjAxsA3xXIn+cFBWsGXDXg+usRhIdcLBTlnK3k1NSzTODqm2kq8ioTskwZx7fMjGmE7asXiZarZ
+uJ6T9Qj/APtLqFBgQ0U+yqKc90pTdqV8Iz/OwIIioVvNQ3DisNm6LGSs+c8MtCG48KwGciuSx/N
+EoT4cxOPMvFQPE4T5AdW3z5UH4bx7QpWZ1hihZ83Pad24wXQGFtzVY2uidbUi7ulrSW/3Vcgo9i
VzVDEgxrGf6xlO94rO0QvZBEeP9oHzAAbDTbqriy1LpQre2fHBqhS615ge39r2AHijOSU2Lc8EXZ
2vPa/UEU53s1lLk5J51AjLei/JQlAs2Mbxnssm5K+dLeQPiqcPLZGUcmTgyxkEM7zuGjOw9pEW3H
8fwXm1c6bpupONI6MnimKjbC6AiykGosi34GXOBywHZn1cQBmw9aviJczGQBgDfSSL/fTtSogHqV
P3TLMIBIQMhNXaRysy1B7CtHDf78nm8/Ix1vvHySwKgjGNT2Q/GBSCLMmCSfMPIsKjvJxFTRGcxq
6qoPSYm8qLpd8PTC86dneSeGcgGygzz0t7LctPcDRJMEG/0w+3Y6j4nAZ0LAQC1oJiEtiRClyqEY
/iIW543PuT8yfn9UX3dQwbLk21fm7GHCEzMezPYtCT8DqM7N8xcJmUaVJwLNFGSi++xWdTa21WRc
tItx1JPaagRNFiVQU7vA1rQ7H2GQmTWU2iWiSss6GByUlmhLJ3xE5phaqTdTnCEs+b9QfYjUG98Y
/DaCqpq9xmBfroD0D+ge+9f3zkRaiIoTPSV0HEo1/GZ0il66Jy0ms+6NVFdTolYJcN5+S95CP4Xn
TA+QAr68qefRSwwGFFSjtNLzVgHmqc/S7zRdVwZCix5iOzXCc3Vv7b029fY+h2GIRQnvbOgGvc1I
hkZL4eU80NmSP2EWm7UMYQPNx79ddJveF1rSi9nkbfjBLeKKt/D9wFWrLxTd6jGpqLUK//ZGvybT
lmX8uETYEqbLCGyHoAnVQsbNXqy20nZLr9vc0zpMqugOfVDuWKqaYuxUasXt1HtzswpFJ4HdZYw5
WsDVzwd4NIXDW848Vb9EbWjI5KptiHX/cTMvjHU4U4vmqUAv3Czqpln02d5Zwc2eiBhbm5G3zkzt
W19hZd/fCdk0WHJBSylqsy6GBQ1cbRKYDlWbfL4VvRIbXvYzYoJOoLgqZesss5/vdBgRKsHfupav
xyho0Dnv
`pragma protect end_protected
