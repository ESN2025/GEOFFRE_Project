��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:�1A��"iOWV��Q����u="�D����/p�*�&�8�W�!�������)��U��e�:�.��u6 �Gd@�^x�5��^�$�lX�K���X��:�y��6��j�ց\�� [�J��?@[~��$oG[�`PaY:�������(�-kw1��|f!�����@O�΍�ߦVP�݈�m��h�:�KKyf�+PИ8��JA5�{%u�����8�2=�!]J�̟�X��;6(�?�ᅿ��(f{�c���	VU��r��K`���&���n�g@���`�Q��6D����,�jW��5��O���\��J��Ø�U���<���ʸ�"�g��[��[�ސy�"ӽ�Fr��y�^c�UGQ�bd:R��IK��z�����J�Hs�4�3D�9xtn)S(�@�g�ַzp����*g����|���k�;ć;�4��� �(��=?x������D���;qeh���;ǖ�.�`��w���E�Q1�r�����cY�����)	�և�	K����<Y'�>�E�i�c\�Vܖ����\;K�i��T��De�08˅ɒ��pcQaa���!e���s�%���:��)�#���8�p�#ٌ�m�3h�	`3��C@}��,����3�×��B���G;�3�l�$����>T����<�[3���܍\1j27�K�[���^rW�E��w�b��K��%m�8�<��	���y�C������vd����Y��]w�&�x�jrc�$�[g�v�YJ\�`U=�"u7G��Fc��ke:B]�1�Lך��\|@C��;}}a@��p$h�1 �3��42��*�%�t������=��C�}�'��I
���غe��"`�a_���7|�w��<�J'��xc��Z#8If��&`҄������dg�BlY=ڱ�ۻǻ�&b]E�&�3wJ߾F���s�G�&f��37+C"�~�S4�ݝ� ��>:�y���������F�L������ϋ���p�=Ά1kR�b�0j��q�^���2sp����/]�ʉjrX���  ��ee �Ԩ��;l �$���ҏ]�xG��o7��iU����L O_4/����DWE_�@(�]�&�����*����u�žd�z�כ�ݧ�Fip�������H���D�	ܘ�x� ��9]79,cl�
��{a���,��10*3�jƦ֣�.&�sq쿎�Jz�����1�I�C�i�Pa.n9`���h�c��lZ*e��� ���+�?Y7�5���J�,ҝ��ڱ��ޞ��d״�zܼ'V��œ"՚կ4zRp2��+�ID�e��p�z�j������$�0}�K>�
�#J���20�R��Vߌ�z�0N�rH&Q�Á�<B�e��0Y���75����Jm�@�i0B���ѿRw����y�	�#J��I�p&�"c���@�,�D��5�����̫�Bn��P
�C,#�����؇/��!�.&��k�X��hh�:����X�1Gw/̠�b]�5�d U�=����A9�k�����i|�w��N?FWmr���K�^
������8�*�cp�x�(�9`�s�����+�9��߭��6���%ǁ+�%֥���kS�b��x;���m�ѿ�b�#]M�[�Ct�i���>,���~�y=\2o�6ϗ�����3G�'�@<d-4���S�Er�8���\�	��Mht�GpǦ��E��Y�H{9�b������K*���)G �2�p��_����y6��_���8침�9��67��R-���sz���@k<��Њ�QxnX������,�)u�"0�x�F�ɜ�%�����=]#���=�E�������C�4r��+��6b��Wn��	Cؽ��JFՔhk�'�U��YM� ����E��F��h��&�<"���#.�v$_����Z����+�oէvE�"2B((��,4�!7�y�?n��{���T=tM(�kD��v�j�����/(���)�٧skS���x�b�2�n�u_߽�rޚc�X�VO.ڔ'�򙟮��n������i���u�>G3E��6FSo�-��f�x�m.f���pAE�"Ge[�+�<�uW!D��yw� ꖳ����/�!�ȸǌ.�l9�`3�ѮM"nzi�Z0��*��v����DN�:r�v�4�iظ����F@�	�P���FN�u V�\0��梆�d/�DB)��L)��1�i��3��]��V&y��z7w��m��h%����
X���^�{��nT¦��	K7ћ<�9sl�k��
^�br�l�yC�)�=�,x})w�I:��>�����u)��M͹�a����3+�ͮ1�pr:n��[�s�;�R� ���/�0p��B�"��8#����I�}MH�jF&�|��j1#@z������I_�MA�Z(��;���ogEM���:7zG�QszF|��.nOO0ϐمk�x<[â2�&���6f�6	e#�WT�� �N1�F'�XD�"$��Qf�-i:��I�\�Z
9���]�\nxÒBD��=��Q	Ŏ,s�-RZ�>�8�X�.�F�[�o��g��h]Dڽ�&��Mn��P �u�k~�&��H�����=_�ԮfJ�o:��0�:�\�� �;	�N���ek��U��'nq�)�8�?�z�yd�W�w�0�<�|�Z�&d�,̯��ᗔ���Ԧ2�U�rE�
Xʬ��3�����W~T�7 �n�JhQ��*U���`�t�$�Rxg\[���J�:��;q4��٥��-I��_��Yr@J[@���1V����ɓ&#��~/��ϚĄk���0ktրXr|���kw}]/fq��I2GO�a�7[�rx�\*d^���E��cNn��$������h�J�]�� �l^Û�������cN��\�����dŦ^�Z[ۉ/*�ْߍ*obzW��C>�,�H<���v�,CE�>��W[�ڙ�+N1�㮠�{+�O 6ݪ!�cL�+4g"E�g�%!���v�c�uf��� [����ʼom��qm�Ǿ_��P����b���<ŵ�7�z39�N�l�l����Elͤg��o�Р�g�V�.J�ߣ]imP)Jm5�!^�3h=|�d`��i�r�|U�������ŉU��j�xW4W��T�_�M��9�2(V N-n{�ζP/��S��1����+N�w��,��4̃�"��IyHr���Xv'�}��&c��P^�y:y-�z8߱
�	��MK��޳@:���J�l����,WĚH7bR���%^�FP�@��,�!��8�v�Q�yI�'㿪�^iHq�(lXb��v%g�.�7T����Z�0Ń>`�:~վve�6(�g�ݺ��HF�{�u==i����w��8bh?��D����o�$ �? �zhBRy�F[Y���B�y�N8���`�5�kQ9럐�r8q3�F�*��RQ��\&��i��@ӄ��n�)�)ws����Q��b;�8��e�Is��eb[c�k�Z(CH�@EjNX���4�L�N���w~)�f�iO^�{��%.���㙷�}��U�����g��[[*��ӣ���}���_ e"�j�ۨ���	ˮ����Dل1)L�t�?��.n�"�����%>ȴ;*@�U��zءA�3} ��p��H��W���uq��s��w�s��/���j��Df��g+�bWg�	]*I1�a�DK�}��S��$�͓]&��[��R��������(+�~ئ�x�l��lW%m2.l����Ĺ$y
AȆ�,��_9��P{�Ƭq�s4�:r���w5bDBq�럟Â��<J!�,Z�F	��X��ą4e('.���R�n�Cq��I���Q=I��pA��P� Yb����'s��oRjB�T׺���㿬V�)f��j%tc�o�m��HI���`>-��* �p�,��4����cE�OD��"�"������y�|�h$d������t\��+��u3Yw��e{p*�hA�m1`��2o|�t_��GD����KWo�,�6��� I�h	&O���i3@#��J2���Wz_�����rz��t�}ն�� �ͦUb��r�A�ul�g��p�)�C��n�Ôb(�O���Gdf�s��'����g8Jd��}R�� h)9�ȗI
�.��T�O��V�)UW�Kه��C���tEH��e�*��������;�Rv��~0��!����(��0�5U��?�QhG��o�������*S&b�=!o�D��|��2����ˮo��W1�f�t��C���0�)���;����Ŷp��W#S%���>rX�)�	j�f�މ����	Z\^U寰"�)��$3o�A�	�{��G���\%� ₾\Y$�6`p=��M
�x�f����\uM|�n���ł�B��v��,����Ѯ/�zZ����{˞C�����<~�L��QJ�9ܨ:ML�߾�z�..-�̆��b;��8	M���Э\��d����8bqr/
�[2L����	br�>�A�s3�)�Nw�d���b����<�����A�;�)�L�w$�n-(S�2�x�@��n�0{��t���u���bk�8����������������W=t1�&ʇm�rM5��
�DZ���h����~a�⨮Ҙ�i臷����åpe�N��~�����K��q�{h��=�BI+X���A�~��_��3Y�Y���~�e��+�k�ߩ���nR���xI�nh���>�M���zUG2NjI
<U~��y7	����i���$ȴ�����
�q��bX8i�	�c��ΝP�*�bH��>?����7���-��}��n(E�ȅHa䁎��vǈ6�k���W��Ok����;����a�0�!Xs��l����H=|k�R�!O�� *)/���76�c�L �:�p<k���t��@�L���X�G� �kb���9�;�*�)I<MP��1�	�c
i�D�0�|B��������(I�6�ʞǡ��UE��h�N����͡��v�����v,��Z+o�qڢ��x�މ>�$�j\gt�|�~��`a>K��].sY�ܑ���~��T�k1�Q��>-�uw67��`Rr�4����"�U�A��!�K�HQ�F>ΈxD�r��`h�s*��=��j��1>p�1���Ume�oi������xVS��%���yj�9�����v{0��#�١&�z`l��U �с>�'hJZ/�?�VI�u�ξ��f�V����&�j�����y��$�Z���a��P�|��܇��թ�]��)냐�X�R�7 �k����Q;9x�\˱�6W&+�r��'�G�È�*�jo}����Nfd�S&�aO�����q|�y�����$�y�c�x��KZH�Y��0���=(�3�M����Pe�Il�9ƶ��^���
�bI���1u�1@!��-�`%ql2n����?V�qC��질w��q��_im�l���(I����WMa/KLh��0uZ%��*Up���>h���5.�&"�>e��Ӭ�c������� wm�Q�+V����7��^�E������ �q8P�-��]���s�-uS�<�7`c{;F)��3ᆦ������%@�����g'7�'g�
)����:`�@#i ���JENޝ���_��[w�x{wY9�!�;*��
��9��
��Z|6Ѕ�M����9ʳ�x���A����U����@��h��W��:���H41Wj��Z��m4"���l�K��\<d�Y��\��98����Z�#�/�!<?��0>o�� Y�?���E�����?3��4�B�B��GQLgomw*�)��6�簢��o�?��Ű��g�`���-�27�Ͷ��J?Xl��a�;O�MV��_�����x'�6�l�[o�$݆	�B1�,@�K"3�"�yֿ��J����K�n.��z#U����㄀���6(r�1,/Ɗ q�� �b��==�-�p)���J0��<��Ō�{���ݏ��8�n����{	Yh5j+#%�-��Y��܃�ŷ��À��h��݇�=s߬��u%���BNɍ�wZ�������������Fd��9f^�����z�t���D�zi?R�E������ �@���nC�h�u�R����_mJ~�:K%�R�T�M#���B��p�����`��w�h�/��4b����W|��Bs���\̈́��W���sN^?q ��I����xl;�6��P?�r�$7U/�Ǯ����.UF�
"C�9��S{upQh��nߘ|�ܲ+��{++Z��eLզ�&]�L��zI3�p;Q��'��SP ���V�$s���[f�c�Z�?�U�F��Qԇgӕs���A{��������^�����[�4�W��I��m�{U�1]z{�&��گdHLJ�"��e�.��U~� ؾ�t(�LS3�s�c�f�WY��)�S��{=0�(a=�ʇ���5'Ǚ��4m� 2�p��f1�r9+7��Y�f�
�'��W�c�I���'�MDه*ÀG�6��s��T�d��z�+@پ�/�$2���k9�֏�J+��;�=E�kt#�Af��E�/��A�jx���A~N��qB�U��>��lYGڡv5���� ږv��|+l��; im�- ��@���Ot�G!\t��ɩ;��h���U��dX.#�k4֙}V�
�ҹ,���@7d�ۃ�V�/��@�ʗaף��,�MY	�D��$����;՟JE����N���R�.��@ձҔ9GW�g:3�U
�2#��9�H.� >�vT_�vkM�������Z+]k��N
�_s��F��c���&M�No^��{�i�$���<�/7��e-lhw�C>�!�v��(X� c�2a�z��v�&aη@ *C;=L��`���q��&��'��1+:�NX�u	�妸m��r�'�)�K�;J&;�@B�{]������<��O����A�����><g_I"�7#�r�WM�<���:?H�>���i�X[qi�e=�ᆟ���q#Ox�Ȅ˫Gj栲�P8�[Ƴ	�MS�ٌ��q	͑*ޭgݿ^G:���
�C�-a,�\�O���	#Ή"=E���d"خ�o1�9QXo�}]��P`�ډ���~_���'%�c�S.�.^�)䖝\my���ßF%�%d l��y�Ƒ��V^,��GZ��-6x���#k�R0�>y��s��)S����w�m|�2�M�L@)q��l����l6��@���F�y똉*�V�u�'��SO�BJ2X�r�A���P�.�>?��s�f��H��,e�b���1X���|((�@?��}��\4����4Ȁ\������U�t���иi~ǏO7X?3J��'_L�u����[l(��2�
S������q��������� �IT�x����ؐ�%��v��-m�bL?�1p*Á5�@c��1���n"�<���k��`�.��.�D��:�Y����B#�SW��ߒ`����Τ�<����� �7T�>.�#F�,ʷcퟝ��'�1�O�Pz<�6n�H�ͼNYC0@�r����F��7���s��UHL����6u��B�� �iђ�n��Ì	]���x&H|6	 }n9�5<���V��r��S�b~�щ��K�ꞌtAv��մ����zko5��Q�{Yƀ���P9���,�I=cZ���Jg�q�錐�i�<%ͅ�����y��	�3�YS^a�X��;�Oǘ)�3:`)�э�Znqk��@Ӱ�J�K��8��.� �S'ӣm�Y����9�tX!�Ĉ�rt���̓>�����SV��(����MN�r�fL�ƒR�$Y�>�8�cM@N��:h�D��?�>���U@�d;XY��6�9�И�i�gQ�;��3�˵�0 i�W��F��S�mV�Ƭ�5o �+�a��9�)[)p~B s)������0xUp��e�!�����Ϡ�q���P�n�Q�x�3�
u� H.���vZ��U=�d*�,��p��] �><��C1��gR�0����8#��Ѧ,_�"�9CЍ��g�ҷj�����d)]�8�8�(�S�m�-t�}���\�Mb�iA]M��^v:�d����S�݁oL^O{�"�L���!�E��9U��m���S����'\3$h��X��,$��:#\�c�Jck_��E<��e3�
҅Z������P�ؼ�`э�{54��٩Ѫ�pz"'R+�	X��tг�󙃄H<���$���N�Z����Qz|����3cΚ��=�q��L���M5�p��p``o�>�� Ӎ ��K�$��Z�:Â2~�aé�2sDd��в)R��n��:��I�*��N)T��I辂qU�ʵZ?Ȁ׉�7�5R.αᳱ�����s1-�)#}go`����r*�0ɦ��/*�a7�6��W��.^w���m4�fp\G\�}ٟybm�ŅDM�'iC!����<�`�+v������Eثb$��&���(�ʛo�\D�9R��W
F'�<�S5&f�3&���Sw.�`E%�0����R,S�;�?(_����k��Ǟ�t�O�"�����i�p\M�/���?íG�8�,�N[�>��ª{U�i����k_���z̓�4�(���H5��U��Z�-
Z:6�#� 
��>4��*��ɽ��d���Oܐ����XA�@'I���R��S���E�CFK�D��m��U�W������7���*��C�e�e6�n:�	+76ܦ�1��fe���Mi�����4֓/2k<~a��DD�ʐOD9��~&��WK�#~@� s��1��*�����mtݪ�h�+5kU#��7��i��5�b���5�~W����ӓ����N����(U�߿D7�/L��6�^\O�7����\6u1s��1o�T ��EƧn4M��1	.Ů�M	�0j�&i��%�d��Wh7�A/g˨�_�T9!��DFO@���vh�w;�N��򟎟���-s�ǿ�U��Pjm
	��OhD6`�~KXW����I;�����eda�}T�}��/�D5�$/��N�\�}3&ٳ���{�p%�ǧ-��z�"e�SvM��m�)�&N����8��
vƯ��v;%�4j ^5*J\��{2�ӥ{x�f� A��>K1�U0���F����yO��~�,c���dP����T���
�6��US�$�U�q����@��=�Ru�H�M6@?�:�'��;���jV�ص}�c=d���n�m�z����㑵�����!�Fd�uߡ-Q�雥���j;��!u�1и|�B�ے>��l!�M!���Od�8�^��b�~S'�����;^��� Y��dKA��9�ơm���d���5![w����%�����>��t9?�$��}�k���O����d1��P�]T^{<3��\>�mH��~� �
�?���zº�~�	�����A]�Y	:�j XZ07B*w���<����n��;8�g��6�*�J�kӨ��ʄ(����c��Ji8e���#��'DuP���/�h���싼�ͤ�>� ���,"�>��/��푵 R�iڿ����i1�ɸ�/շ�\��x��Z��]�.��_$���nq8U���ݕ|���/��ʈ�c��Z%��O�]�$`9�Yc�+ѐ���~��*k��/���D�Ͽ�p�v��g\�^��v�K�Ϩ��~N>�:�|2d���P�K����G�ɢ8��D��Hxd�iU��9�$w�i@���E_�����u�԰�d��B��|�y�
`ddW��&mk6��Vs#��]&�l:���_e�Xt����z��p��Q�ry����*7"*�"��`������b��ׄ��.�G�c?L�C������ayKV?�T���3�7����[����Z�v�z곱��=�a��/~ᅑfL�<���Hۃ�ʽ���޿�{�{����jS�'bt	J^���5Xe�4�~��
��� ���t���V! �t,#HN�؅�)b��=���?�sg�o|+�����ϮΩs�y5��gM��|�c��:#�x�� �sp���ʞ��cR���ǰH�6D�iZ�C.o�F�i����y��w{���Do����F�$�B��+ r��A�2w� 
JLc���}����`�M�d�[t��q�/�Hq���V�I��a��Ҹ���Ə�u:��!צWP�l(h�.���D�R����i��;qLIO��1��fd/�#X.ʏ��8 ���[��w#���J��Lױ �����*��|�U��Up1ޗ
������W
iHO���"�a ���OאVO�y��D��l$D�1�Ml+g?��H��XBENUU��N�W���J�֢�da�Y���e����[t�1͹��=ɘ����U$E�r1ysdx���z���+VF������-#����7�a�M4/<�snc�"��v��&�>Ɉ��#G>Yiӯ[�8L�C$wO}����$���Y�y��{�v}@�pFgL�m�jn'��u~2�����Ul(�ƪ6�|�so�	��༐6o�����%����c�zd9P�+���)��)�ʻ�T\_���1��9�<��^���)mt���E����ˇ|\7�n{�:UAb�n�a�TE�������"�����<�\��9E�7wZ�>& �s�?8#z�E)')ωq�S�e��J���T'�����h���9ؓ;+��bu���[����4P�9&'
��V���<�ņ�y��b�8X=0��}��J�B5�#���6��D��xfK�P
᰾�����
&5Mg �)��p)���?�zJr�XS��F�<-$.��#�b/�L��'N	��#�M�Jt���L?� &	��Ŵ�JP��5< .�������.4	I��~M���>�j'�R�Jq����a oA��͐�ܯ�_�5�^B���� &	�q�#������E�v�F��1e#��N�����Aco�q�\��wF��9�N�/��OW����m���v�>U�p�WB8��tO���3q�YX]���4
{\P6-��cN�l�$�T^j��:S���L�n�
��mW%k&�2v���DS����J7`G4�U�(I�ř	Z���+�9(���B\�><�Kfvgt& _U4�D�_t��gz�,z�t��������D�}{,��2��E��!R�#��,�"5D2�<*�<0������϶if��Omd�n�u��~L4��t��,�!,S�JZ�I��8�#��k|����v
�x76hb�\��zH�^8��@&���)�����������q$\S�ޘ�L<<�R�d�.�v}�փG� ���>��>�L�Z�O��	E,�[G���=u�:�m��`�nm���^�@�Hy(dD�zH��#�0�F*U^آ�X�^�co=dY����?����x辍��!���iX���L���XaLmk��%3�V^�{~y������t��)���8,j3���z��q����
�����
p�� ������k.:b��C���3Fʑ�1H0��i'���4�<��j�ۮ������,� ���*.�t5����A����aU� |� ���!|k�8� 4-�Gs{�ۮ���A
�J+����$�Jl�+&X�ňj���T?
"�ԝJ瓕#	���c�o{<lS��V���KS�-V.h���ꋘW3�ո�^n.W�wU�Y�m�A���-P�nY�aڕ����.Z
-�U�^Ք�1�$�6��/��$�X�� HN��L�Hs�,���m{`(�|��K��z��RȻ�?����˭/�xMkZ\*��$Ҁ�;��T �8�N,_��Lp(.@�~.�Չ��
x ĭ����>�D���V;D����W&�������t�
0�7��aC�m��EG@K���L�s;=m^HE�}�M�Ϣˋn(���^ǧL֨u�zj���-Ѥ���\�B��}����2�E�q�m
���
n���J� �[AҠ� اJJh�F���'�@��@hL�U����x��G��\V��&��\��E�F}|����^�[J�{�Ҫ������W���<�k������}+��$g��������|;��7�у8.�����|��ߺ���#UU��%
��x�D��ww(�ڕ�m+`E�� xT\O �ʗ�~*�+b	Z�k?�/|j�ޡI�{o~都d��a�r�DĦK�@�
����nu�X���"��AC��1X�����cz<z�xS .��S�f��C�/`������1��˓t�����x�#�7������T�*f�c���`"���#b7���(�QL�������g'��2�n�u�*^��dq�;��bU�z���lm��u������cE@YO8g�r����W��m�L�����h6{�}o|~�9�4b�z�61�$)G�t
����Q�N&m�n�9��?�R�J��q�,����1ƾ�@�����s�C{םϗ2/��`�1��]3�D�PC����->�p��b�ۢ�?���b����I)V".������D!���	S���m;-���ʵ�PK+�#6cH��_�+��#��迭����n�j��YZ���쩪�xZ�cS֞(�p���ʩ�W!*�e���6ơ4��?�78s�<F�X��#�Ҵ+�2Y��An_C��G�t��\Z��#�Ԉ�@+�u��o�ʸ����L��Q�O�c�1<§��X����oǱ�;�QG��Q�|�>G��ͅ�G�� %������<Y�7ID���<��o�ރ�o�Md �[P��E���E�+a��:F�l�+�,�n�����(+��b�N�y��̗���V%b
NW|��Gjt�!Z��[E�X�aA�-K+�42[��� �H*Mׯ0���c�Gފ����i_8�����T�.���)�C�[ֻ��E� B��^$�Q��9Pʮ V��<�T�&�W���⇣E%�ob�V�P���HfT(��ۼ��k�&t���уiY�[��t������(�W6�}mJ@�R;2W��AV�fO�[ge��G�v ��G��ϗ�h�(F���Gr ;��v�;d����ąď��^��8��
��*�'#A�����I&� ĸ�n���y�1G�Ŏ�s1o>�l���I��%.�)���I��K�)�=��x#{��_dv��l�$����g�6���}����o���<\Ijr�����n�6|��ֺ�M{���~�[�VF���!I�?,��)o��֮�6sE�w�K��D����Q���׌��`�>p$(��R��@M�Z�C��YQ��?� �+����H%7i�� �x�N�e*S�=F7Զ�x- 廒��++?	j,`���	��|����cvFh��ﬞ+X���1D9��]� (q�#�QB�%�=^)���x�D��x�q�z�x��w��7�CW"9��8�e	)�GG��H��P��v|kV�����S�8\�H�ݛ��6�q��-���\�MDܱ�!+��'�sK5�k!+�\�]�X���<CP
%˔�HKީ�ދA@��I׭h��
աe�g/�����XG��pb�σJ]'�]�{�R��qh��!�AUs�\�?��M��VDEb+�$w��oQ9۴��1B�*�C_ż��rZ+x�J��'垢i�pʻ�K�Z�y����/9
>��1�ncd�ר� ,Q���5+c�f�K�ݟ���;Vi��;?����G�<��[���%��n��}D�ÆB	��G��cѱˡz����Vipwj\T�T}D}
.�Fώ<���i��3���B��Db�|vz{��-q{~N=J���G،�b%Q	��A,��|��'̃
��-�/�z�I�Qr3Z�u͓���^#�\�
�6;Z"�܃�=���4W��K޲���O��k[�羏m{u��n�9�������ö�W�2�]9�)*ڮ�h-GO�vJ��%��Y���9�V�n�ι.
j4��������b(��=9��y��2���T!��p9�Y$�A�BG�y��-D F	,��� jl1�a�x�c��M�^�S��+�|IEH����up2-w]��9'@�b���zl<��A�-ݩe�������_���������-j�a�磟�}���>�xm���2q̖'�i�C�=�#T~Ԣ`K�m �5��g�N�]ڗA#�$@�*U-��C|�R磱��&(=o��f���Z����NZ��'(c���@��5��G��B��iw�Cj>�񅩑YQ�i�[���>�A�������������9jR�~H��N��H���A�6zԲ=�T
<`J�������W]���,n���>J.�>�<f����������0�5�����۟j�����m+�s-��kƱ��mH�ƪ_bkж�o��n�y�ޭ���3�� ��u�v����?%힘�1�H�ɋ91�~ND-��톆}�.#��ہ��e}g}Q���˗��3��`�(�sJ+��˶n������G�T֭���k�.�v_�?��	��l�5M�3�w�OHn�xԝ"{ľ����_��Ƹ���@��	�e	|2�St����&N�����\���j�˘�L�D7�p�yn��~�m.��.ݜ�`?�go�)��B3��v%�p��hR8�|�f��J��9x`|5z���z�r����]�W�fS�L�/�q ��z�T'?d�;'��	���]&��H(�] ��i��u��@��~ ��b`��̦c��$��E��46��)y��,+C��=4��.�������z"w�t�G�裫��j�F��.�b^������!����ڏ�6o�mP��k]$��\6�iz��pz������&�(�}��a|��&��$��O������i~ٿmɀ��̒��^}�yT�COw[P�v ��gl&��?(�\�ԩ��?s��ÖI�I�ږL}�����h��H�A٨�ׁs�q��l�F숫ƇeO����^A�X��j_��X�����t�KSf2�.�5��k�&�C�͟m��n���:4�����|q�U���[u�����I�rzK�?�HE��g>�T^G�� S�P�ǕP���an�Y�@�9+���$�N�ڸ�2?�Ċ�	u}I5w[�=�LrnG��K,ۼ~����.���y$v���E6�cT��r0�q��X���ֆ9��6 <�YmQ��YP�,#�Δ5�h�cb��T�EK_8sJ�i���"� z�,��]�M��e���:�u�����^���%���d�{iCn��E
 j��Se'�gQ�}6t�[j��.�z��o����>̻�w�a
@xt�va�Y;��a!n@���sk���L5gP�t�k�p/ԣk�;Y+!{.R��+�6��c��*�x/[��4;�)@�J��c&�����D�����ʠ���ti[t�7_�V���.И�:4����{��x��.(��Iv�~�Kh�;ഄV�X_���~�~޶#�����Y��bմ��۫z`co! wv'!�\�{Ewز9�Oo�ߋ�6�Oh��C����F��ҥLPzc6��Xq�H��,�d���F��{�x����1J*�V�6��Y�3{I�N�݂���xDm��꟭|�,�^��4�t��f��!����K�n1�[��~o;v�h���0�K��}W��'+�)�{��w��Qơr�v(.��P�:��a2+M�,��ȱh�?���N���z�yrN^W�Qi�ʹ��g�	��en�x��-"�&r�\U�H>�:V�{��]��q�_��� aw^] >[Ѥr��@&gC˙���9#�Bu_O�DHT�>��t�\�Ԡ/�EW2[)���2Hi���v�;@���(_YL��J �K@�,�"��G�N
����=6�ٓ4W���Is�Z�v�?	���.�`�%�ݹaV��1p���s�ќ�����NJ���m�-K����`Xǰ�L�J�Ф���`��ŕ�,k�6�0p,�2�~Tڨ!U�'�}%r�kH�+#�{�w��9�;�8S�kY�*C�Bw?J�m9����v���d����8��3%��~�T��u��&���!9F�=�Yk��8o�N�3f�S;�7Y:�ŝ��	�5G�
�JD�C��OX*�YzLҀ �Ð"���_���Qn��M�K�o��J�V���%`o�x|P���j8�}��y����3��k��<�o5�Bc��#�d^9-��y�!���x.F!ˏ����2�G%�i�u
	,�5�7��D����� ��s��),�/��J`�Rb˯]��$:'��h�N��}[B���G6"�p*��b���Y	n�{$���ܺW�I��2~�^kF�����W{�@mf��I>�ځ.�4jY6�iJ�?N)e�ɪN5�{�C�!���e}R<� Hr�������W��h�Q��m�>\Ww�Oսl9}V�w����{���W���T(?gs��u�:T�b�r��<��d�W �R����n�Q" ��"$�����[�	�eQ���3^i�"Zٟ:���h�W�2�s�����>'���h�A4��1��0��p����8(zTy�E�hÀ�1E@b�YS|��&s����^��@��hIL�^ ٌ'�j�#)B���\��5)�<[pRVćg�(���kW���Xq�1���/TK�3�84?�`StV硞eda���Ihu���d�7�ԱS�G�������t�������4�v��*��� �%5�ʔ��ב�;��3C\8&��r�Ϲח�t�E�Қ�mIH �Fb���74K_�p�4��P��+���|l�4�B�&Ur�q�q=,Ԋ��<(Lz�GkJ\/�BZ���ػ�[a�S]�h�X2[�,���8�=a�@�������N���pR[��9J�u'eZ[l��4)L	i�Z�v�)S���2����J�ٜ=�B����]�?O0�����}��Q�R���X�����g�b�zU&䇍Z��&����;Cc�w�sb|y��&�+d�젏�v��T��@4(x���R��	���EG8����'G�`�}��,���	h?1���~Ag�)�F����N��?�Eߔ|�^XE�� �X���ܲ���&�:G'Uuk]	��W��I���@����[��xۂ`��o�c1鿲�������C�yc�䤖�&����p�aC��Eta��a���gƝ�̜;�w�h��؅S������Ɨ�s�K��\�#��cT�"���Kܨ��i��Aj��XjDB�F�@��q��az�=��wu���V����n�`�c��+� ݳ����W_��xd	=7��J���n���jg����q��-8����pO�Fk<�+��.q{c�Bd0���
�ˍ:,YX��-���J�`�9*�Ե�I�^sӝ�U�^���޼FB �%M�*^��ܾ6���׮��5���e	����7EC��^�nQ��6S!�m<XT�Ě�uԓbI8"H�ӭ��T[O�	��e=�ڡ��n�6G2�W,�_��Vư$���������רeG����󦋞bPM�/�/�i�����)rj�2g[�7?�6����9̑\Z����E}U]	�^��������c�y(���@�� F�kYcvzG��,�9�����K�{}RhH��.��rq�K�сOp$	�/A�c�z�w��aT�0���"_�A�y푪���í%�~V�V�VWy��e�}7NS_�9R�U,Շ�sW���kG��+�ąE�]XҞv=F�����!u���#����+�2Y�����8a��._�F�a��ɢ�̘�g9�>V J��d��b%��$�jr7.6�Z(��a���0p������Db�m�D�&k�ǚ)l���㲄xS��fSޠ�@�8��]���}p���맇{X�.�K�=�c(�3A���0;Z�L��k�@2<���,EELY����"�K�+G��~�y�!T���:��j����A$��8�,X$��fF���-��b���X����f�cf�p�MV��iN� ����V�ui�i~����r7�1'��U�L`�B��|P�����rG��go:>J�)_��P>O�P�n���CˮG*ź(5GE\y����0�P�(�	vQѮ��濳p<PfT��w"Lr�.Z�`����-�q�������fU�6c��Y����J߸��N���f�t�~��:e(�ɽ��*��[��QZ5���V�;�Q_ߎ��o*Fd7�,�ter�e�cL��;fV�ow�(}h��pڪ�zGE?���=f�K�R�E����QN��(�Q��B@ٖ���uŭ�̑�Ru`�\[���徚��O���RD^~��.�J��
�뻟uյihx�S�s��Ә`R�����>}�U��ӵM��S��\x�o�O9�P�vә�8U7�@�`��zh���:DqY�ځ��Y�ń��;��(�9��%S.�1*��ybmO�ZDn��. ���;�g`�#�%�leue㺁b�1 &�ym�LKȇ�!�sfI�V958��B�#�W�@�J0c�p��,״�O���^�V$8E4ϲh�E�l�.��<	��qa�9oe�c}3���r'4���3��޹n�^0`	�<i����~��Y����RDo��i5�rT2.��rs1���Y�N��ߞ$B�lY�.��A��7q�Q�s4��a�c�=�t�K24��Ik>�ؒ�WQ���)�:�Y���:S֒ �Fl�w�+���eSK���4G��/I>��ug¶\��\��~ĉ���{��"��0%M�<�m��_����{cj�{B�]���t��1�t����C�������e�aK� @����h�#k�ZX}D=Ϻ���ш}�a��!�F\bj�@�� ��6u�_�$1j��� *�K8}��}�^�ꩊx�b����C-�0����g-m�Ӷw��:k���OC�s�B�3X�l��׽)q�Y�&c�����8�oFg���Q����o� ��`B+��r=���9X׌��:�)��c��n�ZC�3�<���&������#��1h���1t������b� K�3 ��p�H�
KBh<w-|ELYr���݇ރ@#��D���ޡ}�{eQ�n������5�4Wc�zc�[�FU���Dj��R���̠'دBX�Mp�D�N��N���+�E0y}�?؏�k������:xT��G@�����:���yE�i���&�u��`1�4R�s�_knP,��b�ӈ��(R�u�� ɥ/��,T�+n�H�Jr�'\���ET�ԗ����pD���o��R��Aӵ�X�/}Հ�ڡ�ӌ��J��"ާ���VA���b����xcգ�N�2l�}4��9��U<���Ƕ997U�o[����lR����@���8Fͺ�[i��k���պ�Ɠ��耮���b�E��Y�F4�ÒQO�J�膓ﴙǓ�� ��WY��-�-���n'G�8=r��3��^s"�{���m��OFaƬ�g�y�m&9U��82.}k�[{i,hDx�p�s-����=LMÅ�=(JE����_�\�����6�]{X<��l��#���5~�E�=URG�j�c%�A�����i��X.���M#iCQ,����?ܧ�S��؝�2Z���a���-��*��[���È������
I>p�����+��V�� '�u}XW5�X���ţ�W�'/g
��u���c2�G��f���;�/X�5f�؟�/���"u��`��x��խ���GNo�DSDwAK(W��C)�]��K�+�۵S�R�c%�F�F�|9j���]�`w�-P������'�R��N�x����R"��e���JU�bSܽHrrx_�Vq����]Ch�!@&���-./�~IEB� �ưp<!�C��Vᇄ�@�8�+4�-�Y�P��<�mӦc�;΃�'����7�8��-TX���j��@g�c�ɠ{lO��rt���I�k�3���"�.Ǣ4�Q���M3"�=iNQ���u%xձ�~���{2��9
�����6�U���`���\�����%KUC���O��to5�%��6\����J��[S�z��U/��	��d�A^&�-鞞⚖�]f��F;����*��!���8'*`A�G�s��AP�+@y�K��ܢS�/��;���`��r,M�ST5hn���8FΤ-r�����@��"�H��}	���4��C��D�.�nG�|Q3(`���+_Adx0,D�����u��9u��*��A[p������K�46�(v���$vä��KB-n�N1Tp�T��e��|Y5�NΓ0�l�2ԝ5x���Yl�6�A�A�$,�I(����������d*^m��o=^=���78�	:�UnU�Dc|B�����\[h�Ir;�8�"g!ԠI�1��L��<��MD0~����Z���G�7�n�9�y�l;՚�*�rϻM_��o�n63�ؗZV9f~oOxA�̶0��)!�*���h�/=VU9���џ������9�p��T{5�G,�X���Lb��nxE��3��������eÔ�7N��� �M�����7�n`�DӃ�rB�`\,� o3��	�����K��ʘ�Y5g����ś�G/ Ͷ�B^c"W!��� Ъ4D�ˋ¬�ȗ�f$�31��jÝ�#��y���w�� X��U/ʶ�M����#Gm���r��`��2�	��0��A����7Z����`9���� uo�SD��=w��k����[+q�ٖ�qZ���Lz���K�M�j��@VԳ%����������� ��WSpjE2~�x�eͨ�
uh��
�QeVE`�c�iD�Tk�	n��x�����Uo��)ꑴ��2�҂��W�!7�H蠛ʗ�}�s�C7�E$q��}P��rd�#Hqfw�tJ) `�&���p��"sC{��+ �Hf�m���>�����>1��| ?ۦZ�����˩E$�wb�FKQ�P��4�� ���OsL��	�"�ι\Ii�YU�r=5!��:h'W��!!�z����k�����e^	�{6ˆW�j���(t^������U���R�Y϶lŸ���R@�:ؖ�΂W�V9׬/9R��a���3�J@�5h��ʰ1y&��#���s;N���2N2��O\q�;�la�AHTo_�-�|����s{R[��TL{y��&<�iʝm�������Y-�
��S�x�$���Y��ob�2xɱ3/_t&�LXL�;�B�l9�R@��R�t�x�}%S��ٻ,N3	%��JH��.��PP��s���A�,V9��KQA:�.Q��4V��l�g�]v_�`�R����G�}��P��V"X#���D�;'��|���k�DLK5,�(S3��v���$�Ҳ� �=&i��bɘ>D�Jii�ѐö�S��#�>�Xc}=\C��Ө�윍���] ��8j�:!�>��/l	�e�	��[Y�*�z���nݞ)�ZR5����_b��%lkG/�B9ߟ��dʓ�	 �~���)��@���TA�M���K�U]lwYc�u�3�f��x-L��0y�A��s�5�R�Z���p�B�WWl�ꀜ�]ژԊ�����RneoЌ��R���$Ù�>Vx� ϛb�ܛm�%{��v׬Z���b�<M۩He�D	�_��W@��!�@��:��f�#"���VN<1]��7���D�'YT!J���H:]E�.�Ks�6˖ڭx����@#����o6!>�������T��Sx�`H��0�k��w���@��g��l�sTY�M�'�GQ�����cF2��������t��jԺV��ļ�֧�M����U&�*2�%|, �XD����/1<�R��=?	S○X��?���Z��@�P�'�Z6�U@Ȓ�$T��g�W	�WM���	M><61�6�`����{�ҮǍO���G���:����ǰU=�j��6C�cu;��K?����8r�cͱ�y�Ƀ&48�u�_;,gYe�{��^Q32m4oo���)?��B�AnT�:{�b��'ǫj�z�sXz ����N���IQ���eh�VG���q���Yqi����:����lZ\��}�2�3FS�RK��j_I���G�/mo�7�T�׵|t	 o݂��}�xlM�	�[}Eb_{����*=�F�!}:�6!p/����@�d+�	����[��o[~2�*�$�Ql{n#A�Q\s���ħ������}���:L�b�>�3Ez2]!)ۭ�ɻZ?@ZozN��Ҝ#؇o���IV�/Bpm�P7�E��F#���,���D����)Ӡ�R)߬VC��&���O���/�mxe��h\dM�Pؽ��ӦQ	"����Y���[mO�t�M9��,UV-�� N4#|��Jt���O��\����Zߢp�].{Ṣ�t:+3t�����L��vTE��qg�����+�����_f��>RV�Vo�l�3N)A&��C�����g�y%.�:�4�-=���S���ox��J�2̷�dDJ� |��. �0�s�ya$mC��]��-����DhJ����ÞK��� T#yg�y����֞2�`�z���%��d���9��H�L��E`����p��I�Uo�c�����QkS���R�U[�XX�3���o�g���|a���PԠ��b�N���@g0�[ԕ����!l{�^a�w�۽Oឮt"��6��:�P��h���Zk	:���p0�,*R���Z@LRca�� 	REf�b(��j9�	�5�_^���|y�c�ᓎ"���y#&y�삛I��U��!��_�X~xOވ���*�׿7&t�"���.�/��;��~)k�6��g>�X����� H{��
d#�6�T:|��J�����]ª1�}�����^{E�����z>h넏�5n��F� ��b2Y����̇D��?�J�.3�_�m�-i�(�n��)�c}����x�Ĕ�0d����U��}8z��H�����tc�o�Xһ�����w j����L��f���;B�3��)a�|��У�kC��A�6b]~��'#UX��t\`���j�
�J3_����q����Rh�.�I�T���/�6�l���l�"A�٨(,���岈P �dl-��+���^��%�?Z�𚝧WoL���K��~�<9c��Vr����O�&��A4�� �z J.���i�JZ�ہ�ɶG&�)Gv���בU�f�5���Rtt�4�T��|��"nE��ގ�`��X��4دoի�yn��Ќa`!cox�VN�]uu�u��1���<�ZݸOU��JÅq�@��e��(0���_�x-�O��d�i�|{���d�~E<^� O�A�R,�+��,�6?pЏ�yk��<�����09�+�+B����S	7�#�l~���F�R�\~���#mWk��K;L�M�օ�~��R��k'�����_Og�&�b�Xf���R�4�#qM%�20��W^0���U�9�U}K��ޑs�z ��
���2�纕��{(b������0����]"}���c��L��3&H%���TH�a7�g��3&qڢ����reAz+iߖ=� �c�G�]O������N�P����K���lBX�kd�A�AR]3]&-K�3B�w�3��'R8U�ꫲ0�}Lo��E������@gs(�ۊ')8�?��b���t��[�Y(�w�Pɚ�������_��^\��Wo�)���Z�z�N4��/}����5�'PY�����D$��PXs&�%Ԉ�ȘO�/Ù|65([��C�_�ۆT�:��w��;�'z��S{���-3&k�9�C�qo��DS�HO���OK5�#�w�n;���c<Ҕ1\ �*�J�^��9�(��ܵ�,Ʊ�T�����O���Ӻd� ��y�;����g^B��9a�tQ��+�]���(�MM��O\�\܈x��^2 8��+���6��\��P�=��e�ψT�+�_y����J�֯��a��+_
�u���t�:�O�����w��2��S�����=�nL�h%n�8cѱ��Ua�qs�ŠU�5�5z�A�U��7���Ʋ��VE�������0�%�����k�:ڼ�A�vJ�]筟砦�8[7��4>zS��_�2-����\���ڻ_d�(�i�\�]��I��ʟ�J��¨����fq�u�*��&'�^��`�V{$�*��(�~@>]&�$��t�/�r7=HcjM�,f����5�QL�������t�k9͕{9&+��?����4��Pc�2u"�P{L�>��e�G�:V���0�D��/�O��o�?�OUr@f��W��m�H���ڑ�*ҁZc���3�_3�{��J�w ��.:>o:��
�qު��ɾ���Jh����8��-SU2��h�[U^ݶ�PB�[�wWu��*�fBZ[s��`d5�#�zV (��}R9�z�.�ZQ[̦�� ��
���R��x�=Z��m�f\Y����l���Yʇ����s��xC4�r�;x�F[�h</1:YH���ܯ�oz3i�pW�"1�Hؔ�b�:���
e������ DN(�7�q�d�{E�D���I�e�װFH�e��餸5�`�	�Ȼ�I�|W|r5�"p~_�E�*�ZV������,wm��%��48�#x�����`Y��7fxD��Y/-᭻�sڴ&��t���L#��:7��i�����R�2�=i����$)�@Q;���.z�+Yw�ߢ*�����ioX_��c����N=�|�B ��yW.?-�b��y#?��w�g�&�Q��m�DԜ�V�T�M�x;�;��-VH�n�N>,cr�ӻ�Ò�xk�HลK�m�~A,w493J��Q�J��ï�f���5%K$=^ȞyH�!u'��3#������p5E�����T���v[�EMW=�<%�N��	 q�< ��Qp���F�s:u+�Q�!��l39�$���jð,�$�ݿ+Y*Q3�?SQ��	(�s����X�����xB{�G�%@�Z-IʒE����2G���Oz���Ry�7Y��/��G^0�e�#j�U�Ӛm"��N�n��j�hI�<����I�D��0��$|)�w�t 8Y��׵�$Ŧ�Q_pr�^��KL�TN��2�Y��1�S��P�P�-$c߭+Q����:͓��n�]�7m�L���+w�-�E�d��yc�O�B=Fػ*��j\�L��Ս����s�N��q4/*��q�_�I�pw����2G��!j� w�VOG�ѳ�������U���̉��\'���c�_��`�*v[-�v5�#�l���$�s��.=V��u|���<��ǼP��fyͽ.m�2�
���X������:������K]Z��k8�U�(��ؐ��*��V��"�Gβp�i��5b��7َ��pz��`3 �feV���� ��}�)���g��a�x_�Ԍ��A|��P��[j��m�S���fԵ
h�tA� �=��8q%;S%�ll�N~�=.����J��C��ީ�n���/��s��u�]b�����\�Lh{��ě%۝M�I��*�Sޚ��W]��%���3v=�l��%YN�x�<�����T�TC���`�[m�IU�ݝ�j�rC3;�	CI񁃒������\J��D�F�'M}��k��X�%�Kx�;Ud�`V��ꡣNf�-٘�{�T�K�^A�$n��3�"Ѓ�/t-�D����B4�a�1�^>���Q3̟���6+Z��J@�|2�Y��(�/$Y�|�Dj�	t7�.'�)R��]}�����k_b�|-sɛ�2���-��x'{�u��a��_��ՑܹA�n=�hp�d'~�2�5+~��q�9�/�z����qJL}U��ɯ��A���P_���g"�Q�x)z���6�3=!�ţ��v��������s0<̗z�M����ѧ��\��Dp6���x�_��fL�'0b�HBXYر+�g�8�s�u�F�we9�N�ӟ���g�o(�����.yg�ng/%�G��@Q)p��u��C�:�(��[��Æ�p��hy�M����
c�b#�<���y��
`}
ݎK���*�is��XD\�J�z��b3U����j�H�!�eT�1'ψOv^!����y@�#�bv�=���/LF�b��E�|�=��F�T�9��
�w��ʸ;�3�m��?��H�؜S��b�����~����G�7a�$��"�q~�j>o�s��J�Xӽc�2�+��f��O��&?��s(��3�BU��?����r�Pٵ��?`�U}}
(�Jzg�UޜHOQ@�~!��эF���^�^Z���JHx���P��c>b�!��A�ɞV5�lC=KE���z~G?k7��#�7��i��`�+=Y�ȬiڊP�43��IL*7jnE�^�"��q���6��@����3�P��L���݃vKr��v���̘��L��v���.��0�������H�mV���"X��"k�J�鈶���aa0>s��&�����U�I�!���J�Ub��_�X5ܶ���*C�� ��YY�8��()UlaEb�s~$��~Z�+�(6Pl�vj�!-�A��
����:�0�M�3K�c���|�}@���7f�-������,� W4;q�~7Y��|H��cj�1^�C���Hq�v3�<�K*���ٸ��&�/֨ِ�M�=�ضD�g#��fop���(����y�h��1?	HʗY�>5�Y	l	=MV��X7�K���8#��U���Q�|-D���]��jw�<�N��eO;���nd)�E�	fҞ�X�V���4I�4uu?| ��b����@ЇM'�5s��"�ɵ;������,Ǵ����������[U��p����ś�fL����Y��q�菣�����I�w˅U����;��m�<���Y�u��u�Y�Kx��u��Jd���^s�3f��e'�s>���?>�
<9*���Y9�NZ`5Sj�ʘG�h��נ�<	��$�y8 �j��*�RrNb)��9�C�F@z&�����u����0|��M,���P}��&�<c�D�;�ҹ�	���ʖ�US<����M���HB���@]Ҙh�t���O�v��5o�SH�sn���&�
�fJ ����P㬰\g�(�I��#�aΡ��FD^1NAB�+�>��d�F���:��:��4/�P���~�؝p0\ĥ藃��h�2�1Ko�en��mu&�~b�n�
a����.�v�O��2���i�w�P�����k���t��������2�Ҷ:|�
o�Ӽ�A�~�\�H��u��9�'����4n����u�����;c��hѮN���8� 
��SBl۶jf�!�qK��=����p�E�C;����L����-
��4�QX���t)
1�u�L,KW�Y��RD�������c��GJ� ܬ6}�h-Z1�K�$jO~92w� q�q�]H����1��`��� w�H�i3ܲ�-���S}���e��9L���6o��KS��U("�Hw�m�����(���Ζ&Pb�XQ@�ܼ�`N�����$��������b
;�e�G�{ȃ�N���/��t��7��u*����1�he�Ǹ�vW4�m)	��ڵ�BD��|��	Ӂ>��w�6���˞|#��I�.��9/��B�X.���:쀝B���d<�qa"5n5k����ڂu̨��X $�;q�#��:8������7���͘p<��Ϫ.D�p;jB��ՐU��y���<͗�!�S���[qT��'�9r4���R	1�A�⯭���W���0�h�@�fZ:]jN��!�u7��<=����Iu���)�!5S����F���C8��=;ƃ7���A5���xMv�m��joxB��AAg�^BZ<�����  I�?BkF�f}���i���+�X��qx�zZ���K��<��a��Kx�(;�ޟ� ����xò��4Xa���Q���/Zf��pՒ-,	���wB�<2�D�J�8h�ԧ�F��Iޞx�Y�^�2+G�G��3JI�8�6��$j�Ey�(�M��9H�m�����P�1����FTVXHo�8�ٹZ��n���@>�0��f����m���	CHMTR��Xrj$
����q��'�̀_���@�np\�y/�
~�^۪$|e7ΙxV��f�	CS���e��ǉ�ǃP�F���jD��eo~#�,��J�'�O��b����K�;��m�ee�9�dg�U��Ph֪F\��jD/�x�%f�p��g����z�r����}ϬO5(���z�W©TT��O��x2�m::*��&(�����RT������=�i�8��D�����<���Q�C�rfcI�����p&���/���v�Ht����G0�sT;M���j�`,��@�X��y���J@-�:AR���FeE Ԝn��",>4����5S>RA��䆒l�>�1�݈Y^����ȣ�Jώ  ��`;�^��y���߂w�~<#�,�0w�2�6D��S�>�2R	���I�Lr��D@��@�H��)���98�ri ����1�bҡ.���'��Djv�`O
[��.�-8�����՛P������[�V_�t	��N�h1EI�D��%��b��!�%�d���#q��/�lc#�7/�_�v2��x!���\i{ۘ��KL�=��w�����'
�ڼ���نW�$x��_��%<n.[�;�]EiQ��g�6������m�>�ї�U��<F@'H2%��,����,�h(ֵ��/n�҂d�!
b{�h�iWw�m[�Lk�)y�=��Q�0�E�r���D�Yu/��w�Br���?NS-
�LXЬK<[��{��~Y2�f2Q���f�-@��vR�3u��:��e�y�ȧ�2�<_[2?92�hҫH�$��qWV�s0���ٔ��"H�o,G=�ќ��x�(��	X��	'=�-thD���~`2��b��8NA�=9�H&/�4r����z":]�W��Ŵ��nIr�,�"�
}���
��������"щ,��ܶB|�S���K��u<g|�>���/�7|K��Pπ+E� &�U n�O�$ގ�x1� �!	8�:LИ��:#���rJ��hu��RZ'����=��i���(c
�[.�%�M/O�;�\�~�%�0��X�#nh����Qb�巟\{�
����!WWP��pIv���D��@l�;dc2��thڦ�F����b��Z��d@.�?1Kd��9��؈�.d���H���:������^�a.�3�Q5�8���Z���49�Ƒ��7e��9L$Z�DNx<<0,,�c� ������*3p��#,'����gZ��^Hd�@�ї�>jǱ�2�d�� �4�K#ƄP���1������:H�~��ds,���{1BN�:�b�J���i��4������m�8�>��1&J�R��4[
 �w�h.Zq�g֞�٪���{�Q{/7>�E��kw1��{ l&�dy5�����8hx"#��ꩊ��t����.�'9M��XD+m����F�q���@�f��[&U�`���9���'q4[��XIT�3t�r�8
2i��D�VŜ�*�