��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:'�E�V��?oW�v��/ϩrw��9k�]��ohGL��PԖ�8���`���yAic��b2uB&'+r�V� g� X|z�έ]�7�)S��z3:��Xт��Z��܈�L��i�Ǫ��u���a��m� O�]�u�9�n�/6��S���FI����̻�'�m�#V�6Ł�>�_���l`���,�8�ŧ:#�~k�wu,<wu;]�]��RG�_kG��S�[/ʝ	�̾b5Ģ�Q����4���j� ����r|1����:��[��x��������y�Jw��}a�F�;�݆�	uMF�u*���^���@������iW�?ZׁE���zw-�ff�����;���<� �L�$�F5-4��m�Yד��.����>������N9�g2%<?���]�:�Ў� ��0�N�^���ϸ)��D�8��$�t>���c=� 1z_bF+�@$QL��+P�*A5�$^��T�JD}.Z�����x�{Z�Q�?8�<!�#��
n��)��678i�� T)��$�v�����������7�� /��F�X�d���n�biM�v�]�����)MN��a]@K~!�Zٔ�gM��t%�=:�J�j@�N�76F���Q J��CD�R?��T�y%](�9��&|M��\�e5m�#f�`���uh�Vy��h:�[1���4���~��|��Cw�dH����LE�RbQ˾��K��}���):�1Z�3Z܉���&���yeOʯ.E �o�=��X����6뛠J)�M�r�a�\��zyfg�|���\L�1�o�7�5c�7�`��#(�v�ğOx*�F��)�J�I��s�w�1(�P��Jfw����sRw��
j���ʵ�ܧ�۱�_����H���ߩ�hBE��ŝ�Ὃ�
^l�D��F���y$)���_�?{�G��_�m9�V�BG���y�-38t��J'�]/ˤ֣����`@9c0��Q37�C��:v���z�>�����0�ր�d{/��?�g/�"<�t����n,ޮPO梅��J�\TN�TH�u��*7���GίH�����H��a�@�
ե�w)�6�$Y�5� |1�b�o ����7���9���z��}�zG��'���;��	��s����dk��9��,����!t�f����]Ļ�$�U4�����޿>��B�J������H�f��7�ґ�7�Q`ݞ�сZ.�h�(����*I�!3�����ؔ��?O^>��[��wK_��fbB']�iG�>�NW��U�Q=N�t�.��~Q-�����f��L�si�����3��X��>eA��2���Lu��w�@����1�jѬ�+���$����D��+=ll����p�e���+�� �j&���(mk`?��ޕ���^1�"X���@�t�r�t]2����ER{>G`�Ӥ�.�c�s��~b���*W�|W^~�s+S�wu���$W�Z�~��39�6���Roc�NF`r��WT.��z�}�#�K°���������vP�Bz����@;R�Q�}4�W��'���>�4�	w�����d�N�l��t8�C��3'ޒ/�	�F��5(r 6��N�EƼ!���/�wl�5\���-�9J���=�;�r��v(���ٮJp�%�--��q�g}����ۣ ���x�*Jڛ�ǳݒ�AkQB�����y �������/����x/�s�"H��&�-��I�?%�|԰ŝ~l��ؽ��!d�@"��/�O�!5_Ǯj2�B@йנ=yP1�`�xx=,����	�9���Z��K���1g�lL�4j5���=�����>��n����[4\�:K���c�U�w��<�wg��㖊���Ք<��1(C��<cR?�d3�F�g���9����Ә`�_��g�I�G���N�8Qٕ�����_� ʥ�I� �7p�_F@�B���S�N����8�
��9�?�zpB�
��R�(�0��n���H�lL�ig��Q`�8ߒ�D�dc8^d�؏���1�yV4��C�}���AN�A&�	�p�q�y]�?g������b�U����ٺ�C�}��*g��j�l{3���� ��� R�_Ś^h��$!��9=��3^�`�)��*~0�~9Ɣ3�~�i��H�9��c��ja�3��\O�Z��O����Q�/��V'�i	��0|�lD DZ�ں%m#��:�ȉ��֬��9�>/͟�c�č�dn�<�1�o�"5���D*Z���)�����c@׀�.�/���=�F���^qy�ԃ`�MR���C8Hr��1�ɉH��8��q}� ,B�p@�$����9(|<??��S�J�[׀*�%�9�y<+�MS�'�+���U��0u�))Ô�UW�����,�r�:�Z�^S���/��I��I2�$�+�5D��4��"YV�ΐ��"Z���Uol�w���8��uI�� ��E��q]ɧ�Y�SV�-�6�R�d��%�A>���L; L�Gq�3$���E����䷞aM�Ieڈۺc]��q7,��;���i�s�x͂��[>�+��a:��k�]��%m���Ԥ�B�.7�"kӡ��V�,'p�@ȱ<�ow��?&���X�%!�PG�#.�[�Gt�S��u?F��d4����L���yk�Si�%Y�d ��_�TVK`j|��x=����'��]m��t�����cQVf����	���h��ƃ�w�×t��4-��}�T#I��SO�	��G�J���G��R�8$O�� �j��D���5Q���>�"��Yj�vxz�t��~�«���jU�/��d�_ ���x(��q�ȵ/3v=JeQ�:�����ʹk�㐀 6��ѭPr��fgG�\��0� ��ǅ{;K��imt�Û����(.�vBln��ӻY&�q�?^Q����5156Ч�3^C{?$s	������5�V�>�X��Rhl�DNj)����hM^\�O�[YP��.�p@Ss�.	�L�ȉgXr@$6Y��C�@�:]^�[���v�bé��É�~q}�݆�l�>����x���d�J�#Z����*���B�hk��C �g3\nGv��9�]a���5���hOnb���;��oZ90���y�]P�<����*�2�u�f`���f�Uٯ�"��	�~^�|\�!jf�/V����J��s����!�kR;Y�y�������-�%��#�mp4�~sr�?)�_�ՓP��=��<��%��y��(`Ʒ�{���1Di�B/;(6d^Zٝ�k��ɷ��c�-��'�X��HC�4��!j�{*����ۊ1%_L=���� �j.�2��y�}<QCpC�,״��y/��葊��Z���t�
%1��9��	�����D'�E�S9�:��`�s_�c�����;�V"�غe�Y�(����f���ˆ>�����
|%�������4�˃��$f������QfFK��w����������t���R&���\��X+3�v~�]2s�:�������9M���f�9B��t3+��+�9 �Ă�F�wF���n���=̃n!Q��[� }�;���"=�w� '.�r�j�%_G"_�y�T�?�rDY�f�$� &UX���0z�SĬb�isK<�
��Σ��= �R�3�3�[!4��,�B]̺���yΠ�a��.��>����k��o�m[�EPh�U}t�;����5jw[N�$s��H��`+�����䈅ʺĢ̾_@(����S$#)@q�*�`w\�y�/�W���� �W���n!���4���W���S���PAt���Tw��z�\2�))E�тe��ijy�yۅ�M5�E���),⒵��ta�7����8͡����!1 ��P�a�	�p�����Uq�^�M΃�Į�꟡�J�'DTc*&���h�ڢ��f�L��2�}V]�?U�V2 ���.�XZ���*���L^��:ac��+s�;S��w���1�������TR
�ub~,遛p־��e�%�v�3�/l��5��?�Ͷ�����$�ۋ�37$ԉg�(w�c�ֈx�Q�.�wN/Q²OO���l� �vʎ�[8?5vCR�:����+���.��v#�!��[Q�tKr�����'~�ޡ�����)8�����"*�vzLCh���bt�q�A�f����<u�V�ئ)�8Vzb����S&݄%�9y+N�ѩw�fe�N�1����ˠX3�S���@��4�,��*<���G�2�=n�|�3M޳e�޼k�2��9rt���S>��55��xq�=��,�l�kM��=lzM��� �LJ��v`ZE�r���'���;�,>OHU���ΫG�����b�m7Z'��k7�1tP�81�H`���*�.L�*�*��\t_���/�u���l���iS��3V:�I�fH߯���-����S��!��"$'u�
+`n��d9siՒ{�� �4p��(8�=�{�m��Z�|b��l9���IQEZOZ}�#�D�ڠx�N2��hUr'T�#�RQd���<�z�����<�f=�����*⻖!�
�Ou�A.�@��vW	��(e9�*Ղ���K�Tp�+v�r����ȱn.V��������$�Ї��)��l��ϩRx>wq[gC�0I;��z<��i=�Ԇ�B��=U�M.$M�G�J��i[���3	M�1���|��[�8�Q��p��z7�E(+C�ڊ�J[~����O � K_|%��`ĺ;�%Eh��Q�Eh���>��̮�-�+9�Cg����C�s�������ӝk�T�:�A�@�R6;��+<̍�^�:��J�w��	ߗR�&]=��t1=R���V#��5Αm[r�����jX���)�[,c�ر�v���UO!v����7J��d�uK+L�*���a4=O�>ot���]�ypT���k�K�#����6�&�8�R������F���?�d��X䲠]�43�ݳ�E3㻿w�S-�e�EYt<��
�ө���D�U�V+�R�6�IV�Y��eCZ�d���dR[��-JG^�$p�^��v�2f�I���p�^�_*�l�c4 ���O{zf	�f�nr�c��B��Or������Y13-����Y�l�KI�o�$�[����F�7�����?�1�c@���=uM��zI�|~_"@;S�S��
�j3^`�N����%�e��0���p*�45',_�զ�q��y�'�L���l����%T����ծv�L�t�~W��gc����xV�p,	X<Q�s�c>v�I}%(�Q��Sf�[�%���AKrJ�{�`�&տp
�'�@�b����[0aGF��7 a)XE�\�B���wUjN9�@��4�jd?�c�v��T��T�=س?��9m�
g�fo.�*��*F!,�����۞^/�v#!	΅������+�r��A��"��c�괁�O�9��F�c��bpщѣ�-��K�m�U@��9�'�8ǡ����z��y�ϛ����a:e��\��XA7� 3�O����/?�oĸ�����X����eg<�T����]������-cCŴ�����ڮZ1���vdu �B�� j{ѕ^Q��hN�,(@ X1�$E!l����.��Li�(S2�A����^	}��
4��,����<�.�8�n�7�e�C� �!%�p<���3�
��c�0�/�~	�0J�"�];��!H���
��d��D�Bh6�Ғ=u_���9j���0JMN���;�d��T� C���2�_K�����4 
��?�����3S�v���I���̢��J�����)����9�Ȕ-#��Z�X�� c5��p�GB�������C�� '{�p	3'���6�xs�0mTSez+$��s7}	M��Ņ6J��Jd�L���vA0J�C�:�MV��J	��y��8���Y�ǹ���ڠMg���l�$n �ތ��|��2sZ�QF�EC��\�Ś���S�Ď
�<�W��m𻵻���e}����ݐ<Y���pcm�7�DuV?��,KhM
<��m�!�p���B\���Ƭv-�*���g����t,(h0�C��$�;:�3�[*M�o�~嶐T�K+܈�ޒ�1=�e�ˉr5C>}�Â��VHE�b,�NGݶc��/��=R�����/4�������g�	�.��[jFe�7!D~r�>ϫ�^)�B<cxᖄo�n�`J���!8��iG�@�9�5E���{ε 3��	&:��AAw��&w@�}��p#��SV�h���h������˺p�E|�K�Ie����_�k���@���RK���0*�{lW%�7�6A%��F&@��,�L���pdO��	�WJޞ�`��~� k�����Z�I��i����̿��kT@��7A{�=�q�J�v��>��s �7���	����L��Se�6ʂ(�ni���M��"����GL�\�Zբ��vs+}+H}��}��Dc��)p�E�	��n�u���g�S���������v�]�m��J�#��)s4��y�u^+5����\c<���#F���
�ޙ�Y�M70��0!�|'3ʹ�ї�kլ�)����w�q���j�9L�9���v���RPӓl���X�k����~����ѭ��+_{�{ ���L��s�|4J�dͮX�S�y�K21�П:=φ��p��{X�VcP��[uy����o#p��s{	Q�~�O�I?�gH�,�H����,#G�įb�2�jG�^�W�-`��!ȝ^�V7RtE�@��UV��ܝO*	P�UG;�F���Q��ч?�Ϝ6��48���GF�bv��$���N!#�lmW�J�3}�����'��m��Y��%�3�r�ؙ��w��Þ�K�t��7�f��bf�1*�r����X��ʖt!�z�c(-J%g����^fpN����H��	��-��mT\& �"Ii�6ȵUpk��3} ���:�w>�R*bw�����ؗ���6����