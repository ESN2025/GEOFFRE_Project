// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ouTCQ6Iqf07JTcpS3CE7xiDQpBuGbmUStD833w3PCAy2jh/AaOxqDN5lf/LvmlyuhAgC93DCNZ3q
mnl8RrMaN3vFUWXf73a97q1N/WJxXqQ09oSEnRHigNbvn/NhZ/JlhlBuhV3mWQaBkT5epNn2F353
S3pwm+KiaVXNie0cy5bjwPeROSeuuygoxtWYxS5iQioeukrhM4p1pDo2UH6hPniYWVme8t3qVlsj
7hxNWR+ydINXiSaoRqKTRvfchmbCzyWinGpzqYWjPv4CO2Q0lipSSIdMNQapox6jdKYlVpdhkq7K
mZNEXv9YRxh9mwv0qtJM/ddDVigFoAYeQ8D0bA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 12880)
/Fd8HDQ0myRaYW5wrTFuH7sZyBcs05zLkIJ39uwRq5lp0pxqc671HvqVE3ZNn2+LYDLDTVaYoKQq
n7Je6W8HAmagpm9TukuQ9bIP0uV5Ro7Q0UpJobx3CXz6Mjpje05c+tQz7cOd4mVav6voIbiJoLdH
xTe8cR/Pq2MWSvgV3I1LQM6oy2B6H6+xeHDX/A9XtF7Zg0UwxZVXAj/sA7jLO5LMFR9bNJMW9wDW
hsvWRk0/L9W0DjX5QeAU9wz2AR61TSAhb/Uj+HQgL/L8k4+/+YVuBjxcwcC75faczhH38023u+5D
beP8RdSVpDqSWllRbnGtdFEjOgxcc9xP+aFYb6o0EOF5ds4s5tOEi2TX6plA4nYzUAHbxemw7UHl
Xif8jxsA3FyfpWfeDxR2ZdSPDwKPlsNzEVqEFTd6zmly5rbLPdk6zm7YdRBk8rls3BQ6GlKMIKhF
/pNJKkB7uQXqIxNwWMp7l7PHlWYS6eqStUjLzHvqeL4T2trpDLxqxOfsGPgYaTTZhUWycVj3YCPp
oWU0p2GHkORbSCn7JSBShyglPDZ0Pfej0YjF7in5JnSHfR1J+YnBHPnq02ujdX7QDXLupojnjZQC
euSJTfmNi+JhjDnQOmc6BS/HYgoHKMwgHqX2K1gwQMzdGXIAe8E2s4Coz7orlOe0W6Pp4pCiFYbg
Xcurro+MH5sSqYaCph43uvOYhIbG90dTNaN20zfB1Zc7qrqH0AOErpVZdd1M7wFukfg4+XXpww7+
qMoiInfhAz8db++1QvfYbsHYVQP0L3s16rvifmDXfwPakgMBInQGQ8zQO2xcd7d/3bNHxaFy+Rsm
ZuSFgnaP/9VFUjnMEnk9eieg2vN+vQtepD7Ntr3hBAn7n9zKMp5j9u+TLRuBnbEgaCunI367RQKc
x4ayryCsAq9kmlYSCYXwK/hF3WYsG8S+Izsvb6fzN/BSJsTifz+gH96ZavM5zvUdvT6I5GRw9dz9
BMpV0ilhA1v5pqOng+7Svn70c5Oetn0qAIxmv5f4fpWD0UoWsSBGE0AbNeqktHhkzxfBwrxRo6yp
3xaxsY81YeBFbl2D6kAT3iG7B36HMmpZ9j0lFe4x7B57NOXj6rSuoi9xqjWHpeOJadXJvcaystHj
1hjb+xgtFSaZGcNb00CjLl6r82y5S6htw5c3O89y1CPBuJXVtVvoFZp8NNWgt5Pi4YBmuP06HXvq
cTW4TM8b3ID4F6pmtrHE+MQYtNnHwfihQy7xmaHT6kvrNhNP0fqNtKlmxVOEkRKHxT6sVfRHkJyL
aiXG6mn6TTmo40l5xBxLvql9X8br8eCukKUM/pWfhLJmUukXH1dg8t3q4iLSEbDkYXKF32jTbwuz
bZ5gc/kEJ8g1qHp40CWfOzXmUcJGraTYIP7plB6w0Ti8ln+rufhBTNz04s+brbuDJG5T/zsbskeC
aNTwPF1woJxZG6siLlc05UHNXt1bzS7KX3NvBizO20XCOJ4BTEYZAQwJqJiHZFYR9wpR1P1vuXTB
p6yXqwpaqlYmvUf2sKMM69szr+1CayDP6n9ZTPShSdEWv54rgF57VK1APKzyjBlGrN+ARwg2d+iM
uUvhnSox3z2U92ln9qoyho3g3FwvAwzEXBzSre4JIyTqyNeq/szDGp2jrMtOQbmnk7R0QbLCAAg5
XdiO6tMlP3/3bMCbEmQoyTJjeMKSkcHaMzsXvQrpKDuZO4kWmT5nY77CrR55HjDYxf5uWB3s/kUk
SzGkhph/p+JBOQzBq79mavOdO2jKvex5LtPdfklVVq+HlpI6//rMQZyNWwKDMg7y4ATHH8yHXuus
WPA1NV+G1JAoiLcofvHnGm26JS0leLTPuQTLZ7l38VviVE5hSu6/H4nGSycS0qKPN+wIIENjPH2Q
xfXo43bWZzmRyadzWTv4j3AOr04HCBwXSZT/st6H7NF0LCSd1KjxDkgnFq19MY70lNirYgFzfKSt
VovvgTGDX05dVfOiB/kcBLqL1IhsB2DZYpchSR7ZitYoRSEfGyeQFMsnjVp2kj+d58Crai/T/pCZ
wLdFmGluY/R8pnGGenVbw1a/U/AaevAh0D93OwhGgG+XA43G7emvsmgucwApFjXE8fiRL/1x5tkS
PcdQLeZQbq3g46+nGRY8Rm23qxAfVjJy8OUuaAKJwqQt5g2i8LhW7eyIYKYwDdzrAt9O3xVj6ZH+
4aQ1y2cxGfCOJJQtwHhvQJkurDpSPRe4MzaNFhS62D/ZvDeEs6LHdZahZTsDieIbYmc1VTc1S0U0
2Uzulx5ul/X9ccVUJpHP2vULZ4gUvbs7Ewc/6c5CYpUF8e9szbgO/7EptJ6fEy9/XhArOz60+172
1B5/YOtYcorxtIU2M+av/2UmnVLdKXkIT2mAzaprD1bwHG7yRahJ2lzfEc1ky+jUZnEmhl4QN6GO
fFT4Fvb9qzeJgcAwqmhBrUSKCQnm8lNMhm7ZvK3EzqmVPiSH4IQ8+UOl5UCWOYgcqng6vbFDvT/U
2y6vxLTD+UtsA3r7BW6PRdR+KrfMXtV/KhJw0tJ6hh+WvOrYFIdAjAVVAZEFXYl3ScMixbQDo5lU
O6ljj/nig+dbpQQRczpG9DfUzeNtl42JmJK2AtaPrBg2X6ncziwckwreeRcC7sGgtn3xh0uEO5VY
yLIYdu7cPG366/4iUZT0O09EEkscYP0b70j8ozb4hHqlRnXRkzggEreAuUK7ybOiaN0QF2nI7U6F
yblCPj/d+XgGTtsXqaMGKVrpB7AhFPCR4tPdmwW09wJ8rgjjwNtmnnOd2h2+VlwdTlgnt7HmhKuv
cgCGE8vacHyzVfsTaTIaMgKm+GDtd9WpNYrwKHRNpA6aQjEcs7QUXSSl6cHOWi5685wbFOSQClOD
M0c1v7O437nguK8XU/EkyVzyqiiU6/q1zJyQ1aN+qOB+1Zqd/UBBcWHMOvnrHXsqKNflqKoR3GrC
HIe0oSLa5CqwAQXZN4nlmV+uP/gWj1bu2YH8wTxgHeL7QDuYtkDxKfbVYuJ6A8okmqpKkN7DRy5q
TfIgHENsIhiuI+JJS1DKYqzQVN9SGRG4sdd1IGjU1Rxm4rnERnvGj1oaY07JFOVZweD98H4LCFyT
EIB/ML/Q3nGaDeg+GThYRbnKsb7+uof1wOt/FDrdkpuqHza1SQAFWOkRoiF15LHKEAmonm9YBeKI
a3G+64iYOSZo7hML75gq1qkyp9LN3D44DOhjG85IExX0ais7VCcewaKS3JKW1te2+mc0lVJmsnhG
eS/jaU7O36ICkpfVCUNHW2jBFGDrRdlevc7+sqTmq95TR6o4tQlS8uAGXe/zbz2LwqHA1w1wfth7
cJd7+jDwcx3IfYdTcqogIfqZr/jwSwxR1xAN/o+wl+GjHqXbbu9Ajt3FqPCJ28rFhTFGhuamqGCy
MO31krU5Gb8HoFwRRlXIvgUhwdBWSAyGkqk5DF+qqhfR6uPCxfljKCxDw+A4NVtlfjwKsItMeKhZ
ll9+m0b6O5e43qWYrQ6b/wFn9dogl2P4TxOhTq6zdwucOBqYepu4IvxqciKXWX/DU2YfMgyLoDNh
ICBYeEBEKLjxR8CJzndaSE0OPfuSFmfdatcFKajKZhI4Zz06i7QYHQWraBCqjhRCUZZjBxcn1guG
dfQ+Ei4usOEHmR1M+3k1N6rS30myO23WHklN5MI+suGh42fxcFDw8pPZxzQ/rHdRgbSqYIM8q/y9
9jUejVYapF9iLZ3qK1/AjNWEhbl75d8Y1i/w7i0F8LqQznC2RFyehBPPCIk4jRvJEpjg5mwILAIJ
lUxZL76nJlnUaGH4mzXmrH70d29l3lzOXgFPf5G0iwaRWYfjTB5wiMcPFwypvP8/0VBQDxSf5anF
Qr7NQdT81srNHXg8td3UwKN4y9jIjXbU5yE4M0EgbU9n5T+6M4dEkSYVwYiXBaYI1MTCRvvzV/mR
Db4RFeMZVw64BssY6N0F6qf4+H1q803DhkkNHPvMG4ZLKcQriXjvkMsScIrlUbDlX8yJ9tmxdGjy
qkiuiNHn34bHdPH6HOh7zHe44SYAEC/kRl5WO55rzhSHJE0kDZxgbKf7dEOuP0YcECfEFozMrrdO
RjSouQVAkpZqrzI4LaMf9ZdgNRsj4w7fGrL7d54asiyPVC6b/Cf+/pRX7UUOi1++DLQtzLjdSUiT
ejtbW6XYEYXkq1C7N5bpK01F0oklKuFHkrLXKK1g1Yvmal5fiNgza0AWGcgTU+J1Y4FllwAvd0E4
Po0nx83W0rR8qnWtPspki/x406iZlLClwSbSX7ziGVn4TV7ZmOGnk9U4hGUrmb28D4w0cEC0IoKE
4DTulhFyVgzNzWDh3yxfy6xJINp2fSBfSMKHXRJfBhV6PiszIING1zVblmFUa1GEtY0NfczCErYx
QjROIZNOrirpV/X95RBq6KELtAx1zhNAt9hh+elf1gSP6hAX7APiLj4atnGfSGVLrBesVZ5qi9YA
tQR36W1ETOAx4UKIFIQOdAsqrAodZ+/7CQiiwDDkzas7/yHlH+obApX4GYpbOQeqwkaWhEkWRR5r
bUxH6GZLl/rhq1VgQfavriuV4VhYAq/WJBrv4einUuN7ASAe3HDBcCqT1jutyrQqgp6/bDeHoKT6
g+8qpCRIqJQ3B5ZHkWMe+V1uqOZ7QjIaqmXm/KnfH9H8A94kM6Wu/2zuQyyVmhMmbHHCDaU+F3Ge
LKJSYPR1svRsO6nxGCY2HQSsjq0jPbl/LutgWpcn7hX/0oIOdg6os9MzjQ7beOjRpDKkABSRftLz
bOxDWA8vQf4ISzQlzOh1+WCpWj28hsKKSahEeVHCjJtqAYase4gDFGy5VEhz+E4eQ2bATzaHgQUH
LFFkCwWzpSz9WiJacUe7SUIxNbo7epGMlR3ZB++SJ7B3nNNC6H2+PF0hyXac1v3RuHiWplCgL+Ls
tGC1KKviq8oJh/UaBCHdOiHxB/Ys7edfEcFzHbTFBQhcZTjUex2RRYU3jokVCpTct+U2j2QIjWRi
c66BZeRKFLN7gcTbWIzlZpk81db1so4YIh8Ta+uEMX4Njv1tGuhkIgch7lk9Qj6nnu7uws967foN
RaX/F5nStzpW2XFeICv6GfwFdo3DJGbK0+DDTnOgchvqMgFpemU5Mh0BxuAuFqhci4AyzNQFWe3s
wvaiLPmGYFW/SAVH9jjfe40Ebosz53nautYkkX5SHBj7cj7BodCWDMjHVZQ88QHD3QtxML0UoOpC
g2IAeG7xhQjeZkwkkAD6dEJZcTaGQ2ZyWtL0NPGl5imigLWSJZ3N4cHSABejaXjpCnQW684bVW+t
SBL7HEqaPxFNJXhQ5xSNoy9eCXA4B7+WOlivIOZT2VRg0W5UJp3n/HnZ0uUqoJmGyF22KwNXVrpp
41HXQFK6I3rItMUeYF+0RjQd/sPzS7FAWz4qFOnxGCLLKkXyHdE8OPe0fMI4h+PjIV/HNuiUkXgy
l2quOnO+qI1FV39C7ffnD/U+TE/KYs4CwfW9QK02Ly+7W8X1rS3Qx7TB7tMrtHWdTSVwqSW+le1l
kJ/mZSiOWhCcRvpIeZQghwF5622b3F51dABvIn/Kz6glQ18XA089eEAPM3XqHq7CUZMl4x12jmqZ
0gUzOBTlgE74+J8LG+Kr5s+56/Yz2ZRRQPjpaHYvjodhVhzc7uOn2V8Fdb/dFf+SY3pTB9zuS78w
z59xYI5joRvJIjHW85buvZG8oYakA2GntRXkW4gj32LR0Qa2J5gU5Ws03SemfcHl6ZLvNhFjWRfK
jANJzsvrycEG7kc/BakIBEJatW83DpQdkhgU/3nLP4me5gyMiTgVSh5gAmqTeEhDDce/+TiQoFTL
i+ccOTFh2c9I+dBLgrEiLaefsCVD3AZImaHPZfMPRIo+gdk76OWJzd1ivyNpVWmUM4Y7i9tf6q0A
5PZTDjM7/4Yb9/0D2uHB1SK8MiwdsurWT7oC/JmZYOeLGKiRf7tEvHLBJjRdCe3N0WFCGSA7i1UK
2h13Lw2VBMSmfksGgk6ECtPz5XmxMobgevOm7SjVfZy4y6y3zDzwfxtmYMSux3nFuDilO1Ek+qtG
IMqJqqHeTIbYJPfrEOrPbOIMWhJo/2UOdDTzypBVsQ0bw7NB+QEY2A6omb3FNcKQYsrTzi9/d3FY
+NzyFjUeo6r3CI3TPqOEjwxoUkERLJnBtd9NLmqakL9601ulwYds7Da7ggTZOln7jYUQ2H/0XRoG
wQUHe1UHZSr/9YJBWtDqwV9oKepXFr+IIhdJl1hBQKqqQgu9jA9trk54QXLX/jrdcxWZKKCsjaKp
Izr2wrBZ/v4NqcsLVIXGUKGfI8/ZacR/sTdylY8tsOiYqn7YSMg3MfrGZhd4ur4j9xGfIcy3B9dx
OlxPatEqWE+Hww5V6/5ih5FOpaLZEbDLvTzbW2ENiHEUyJU6/kkbd8Whp5GoGdocyVc4X6iZKMvX
9tnyvW5KW+Oj7xFSEmZAkVQif5NbsbMgDD/cpJaF6pPFoVOJl6JaWS8c17oTqwLbZVINXpZuTdI+
ckWJEXj6DZhew548RbRhiwOuwTd8dlGfQ46OZjhuMrLe4LocuxFXVilWNcMzVdgIvtoUHikJtJP/
kfWdFyijLURXgZqO2zWG23382DyBAnPL+jmI51ARm4ms0sjmbnJ8Y7bfvfjujiX3/qZl2t9UgjI/
/V4wzLqgSoIXsTdE2CzW1F/NCTqPa4YiL7p5R0WuzTXnQNV21XXD/ejT3t8qFscEF73+OLQ56DFl
je/SL9pUdJNtBMlrFaF5eC8BlY3/kj0+lgXcYkmEf1geuOoh3HyYv62dbX67XanLJO/L/EklXfRt
AK8ZqS37ufTBg4W0KhmZhExE4MkOHlkeJYhkaPWSxAZ4BGkiXAvtT1wwc78lcZcwB5/M/Oocn6ES
NGUt0rODyiEOIAB6rkj/ak3zioCVZezFUN7G98uj6O9Yhkwy0OMS7Z5ynP7i3ZFr26xSLW2wYfm6
EgSizu8SQFMl0fSIADXfQILTR5L4QfpPD2aiO0Fx5RlP1Oh2WdjrQcb/tpEp4mDdG3MqUOP8fcRk
/QEZQhpfTqRwzQDthG74N2TvrMWcG6IiQFIrWcPLTYpXExm5B3eKf5XHR/smgU3bIc8qQK5uBTVO
u2f7NPd+OcCKQt/hL3oDEpzcDTgnj09nQuMSIhRViJj0uVm41W3BF/RdxFTZevuMJx56J5S5/+6g
pXfvTf1mzhcy0rk+hfq3IAnpdaxRC/+EIDV24Vp9vWsBdIj3XRTuafvbOGlSD2s1rmysFNXw78r7
Urdtg4v+OYomHupw7l1gDFzQx/A1BYHOgfdH/6C5b4e2gWL+Gdk6IzKDSD/Fb1UVedEi5GhiiCFc
iBIn23Lt0I4EsZLXT1BU0lKP/hojmUfWyxFa9UQ+Wo3ZY28LiRG4PN3BZjj2gwClLeZ/ZNSc6/Bs
ZM2Qz3sQTXSO+etXUwGpOQazE4qbxJu9PhzhdXTdhilqHPGne/5fY4sHYFij1FgqbiF8qJOQ8iyW
HnoVQpXdi9GzqZ7hqa6b2QLeWShsGl/OvsAeGVIEbdQJGfIpOcW9bIMXEDzRzrapputGwie1QyC9
QY5abP5MFd/UM1fHWHSLzMBzxXSero+aVIWZ8F6jw2N8jrw5P/pt4L5iHZx96oCOR+gvLu/IhraO
/jyVUb0z6fghTIFPBQXLWLKMErhxt4mEmUequRHhcJ86lXizy85M57KtsoOkXfzxyiKv+p/HxNe5
59FkO1vJUnGWsAEXHuiWMqevVW6e+pjRAyg1ikxcHOKo+OezQKdzZnQhku6PI3yCGa+YYsEEPRTd
oPRNJqfvr6StsjyKUeK2RTYW2rlQ8KmgrIJAiJB+kQcBC2OVw3foFhFrP8ZywC1lvpxAYRl6mLKl
ZpSzXBSczqQDXByg3EGwA4uoADAxeR3vT8JLa7ckpuBWarWytujutP52zw3tyWQ/XIU6+P4DcaMQ
3PFjIlN2/6zT/g4pA+c4sxV7g9YIm+6Uahg4wD+mNVfsDZztCp7/Aw03qOdWeY1tM7ctZ5cyQPIK
65FAdMH/lpxOsPLKccyq+pAmKUH0wJbwpS2fr7h9riy7H0k9AGUniIhNjtslRyQ6Rn9L8evsbJ+n
tDiqwdEQ3m3/hX4XgbLsvyfOZF6v3378AOcdkbTnjubGAis/RlSqhH0q3XCUqP2o3qv3P+izSivj
MbvrgPQdHeQPRxhtMEkZVmOl7t3XukXUvW0klWlYQBv7qPNmfSyzypCltfffAnTE8MHrIT6RqoHI
iF+V13p79hLV+hqH4oSAdVLOpOCeCcLOf/zJBcNMGpSp1wYJHgDmvoLq4hxvgU8XqpvMZ2w1vkc+
Ueo89A7h+XKZlb3LyatkshfDOeG0FIOWwWUD9KIIIWjFVWkY+qtQuseeH7Gvy9PzxLaRUi6YaU7I
dMZHN097emerh4TRuGbz/To7WScTOYE6kVuycqWncKGySsosTERGlLNLe6Xr7FEWw+UvSNwRglf+
pH0oGCKjvYufURDRPjeuDvhSdrUCHPWHCOqoX7ls5iraJJW1RX2+/kXsxgiboW/wIEOT4EMkV2N0
9iACHiUE5rSeVAZ/9vjIGAAOyepN4Gy52HMU/8JPJYRuIzeZa2utMqJ8R7DoOFaWLvXx/kaBlL7J
Dr1R2lwGmQ5SbjLFRlB731n2ZW7sLtENcDQXIZdsukYS9C0WHgx43wM1H1sGUbIfxDh5Y+RcWeEe
qjDBZBbCJd8cIhgvGEF3r4D6E5FPn7ezB4rNoDGnFbg+ZJMqxJFHEeYUygXtCTkbbwIaIZJ0UIdZ
11P1ndupQyhV02NPcCa9bXZ2zTy0fsliRJtokSG2JwQIsShzIgBypdRoOuyunhMVzqh6uwktCshP
29VmTNov/WI9BxLwuMsAIEmrh85EW4M7M+sIKq0IJQ3MiLFywgDhlfR1UIccsyi8HuyyPskFenvC
4pv7qOXkPtZLJ/YVYXSRXc01CnpN9vx/5UkJt9QsTJcN1sFnFjd7L4g7Zw8fCSpzTPXViVaQJd1K
C9M+a7uZ7sfzm0vDldwALiFabGfzHfCMRTeUw8KatHjvaMCatyMQt0oON608kC1HVsFahJh8TFrW
PKSIi5Il6QDQpGOrIk14P2Uzow4EvLzRLciFdu7muGkT+rIGJpKJ0Lb3jtf/A78lHDuJSivOU9ah
ojsoEM2RtKp3xSfn9gArAXM/aKl/BLGMvSJj43C8oXmZDbSDdzS+a+mso0ZlMwImvDBDrfvHwwF6
vRW9TqHcuIn6xaKTYNerOQH5N4iV4rHp8fepTNwRlYDB5qFUaglMhd1R6lPVkfBlALIlfZ/TJCg8
23pyhq7HsPU/DL18v93yWnwQAFqT5uWrmeQoI9eDOcQMmGqo0+eB8hXsxLt/aiVDLxzwrYF3QKBE
PNC93qZN0SyGuiNAKARruOon0X44luUTC+7cptbFBzdPDjg+2+vOnulxiLLJZagyG3QDSSlptW3K
IWgnQQYRjHX+5u+EA4ZZb6oOQIMHXgRpbVrfKqCSAyUDoy9DMx+OYk0uMvrZ7UPV11VPWexOraNC
gqM+D7QAdtS337V4fkwISCkjTlGnBUqHzYzlNfSgg1tusOmX4/74+lOOqScFv6zQSBVnp/zMHq1o
nUV4ZWjKd0eeh7Mgu8NOd3g4Tth/aFdXcZksKJplrW9TJo58nCAfeui1ar+5iHqc1XVd0QrEBy5V
Zo9StIcLa+srxxSSC/opgoJ6P+Lqd7cWG/pZRGr3zIw86+Q7HeNx0DLGlKexNBSY438ldswJYg4y
i2DIFcP38eqodBpheHp9n6fKfgGyTbxvQ3THrbi+jw9G4azcQKO2JlQc4D1rjsOJrWice0XQ7dun
+Xi+g3e7/ziJdQ1VVEqVsrunroW9gbgkZXERrmd2x/ZUD0Va36GAxuYvjmoJXLwOlEhWJo4eRWAx
Ud/ngVOjG4BdPvzPcX5NmaSUsGXbl3++hDfa2bDPf/AMAU0BDPoOZSEYOBnPyzCGWT5Zg1QDqb/4
FNZCfa264CoEtCrG5/3FJj8Qa6YpGLDEyaX4eeFUO4Ou3E+41FRnovHt2may6Wx7NCjXtE5Efe4j
zXXS5XMyLG3Ff9H687xe16s6qu/ONiBD1L5o4h+gO/wzw7Fp+p8xaSPB5XQLhMZFidYuyh37vvMl
LzvHj2HiqeUXw+pGBnHY50XxLFK4fCWj0E5XsTrR0VIaxPeBjCLwbPXc50F+WhX2UeZUqS+H5lYM
rkb2PIWhPnVreQZNptJKWZQDhWR1jL/iMIQI9YZbj5/QDJnBFyD5So17QRlgh3tYL4kD7TkUqbDI
xu7vw4m/JDJkMJQgU9o7Y+zOpzMtBvrTIgXTmnlT6PW8WHbea5E/cvHeHPdTQK+/P+J3LOzmY+vH
r8BoHaUZH8Ths6zS+GuqfsS/tTnCbQKdXij11NzVDUa4sCgFc9vZqQy9CbEU4Z56vuIZQwNV9OMt
GBxfnrfxexTCOvixQVwgk1iaWSbyLljuktOpFhz7TFUJ0q9X0OBQ9o7zfCTMaypZiTxBmQWEKTMe
6LpneY9Ig9KYhpa1ZIbMLUP/5AzyLpTUj9jsN6wtpGMSXNZ143k+IdvCe17kiQxW6nbH/q03NJRl
tljzMwcQ0dUCPx26TfME7LxUwHxvuwFayINZuiJIr6vcH+m1cLQAUCC9BWzBiP9r55O6BSweT66G
Om8UfsAMYTsyrqTPVFZOJ59+TP+qMpJtTGz4eOSO6CyX4Q1kYWyQ7nVBX8U0XBd4L81/Oq0eSR6z
eaXG7CeJpNbqUWQUUdWmCE+wAFVd7xtCyihLkw8XH6Ipuw0RZIuWgRli/Y1LyWzzb6nDHu7l5BvZ
W0qkaxe3nl8jrEd19GXWhfHPm4Rtab1sNLftGHVWJ6ZM0r+VSDFAVULC8st0ruScprvuBlUEynQk
Apuf5CLUhpGtU03n5LyH8BeXEy7rkLT30CEKiK4K7TqYBUCKsB7bqILGhnB895r+BQCrzRNVvcOj
f1NdEkGaedlZ92U4qEvetPkfI5BH8H/zbtiBsgiyvEElE/v3o7zwuIbR1w6YGz59qmpiwoHUKmoS
IdHo3oCMB7YVBIithPPIGEbP1l8EdV1aUi3+EVJ4Nb5x8iwSBjKzuuaCI3UBY+ouQuloW0OWKkM4
AjU8D4zCjII/hXNS/Sxx0rereShHatlkdyaoN58e/VK6O7nsqC/tiLoZ+EQ4BZmpAR51861T5dOC
oP4wP/kXUc2CL5jjmT0NjoEEC4YLCuq8WMqEn47XjlajXnK2wVhwonBwSlIw3ymvORO0j35NgT6G
a/AYM6bn+nO8Dt0vjseoireWAa8wizRoCBdhvhM3dNgDMNxW4JfzGBHJj+16zlfFM+rEUnCYSjIj
66kLYb3awdQ9BQPTnRQCoPbn29E83ihfkd4Z1Qa/bSo5akByO8S+qKEOuee5n3rJGf3jY/ZH1WY0
dcqIGIacH2dqndEfhnseimVu47+MlZpql4m4LT/TjFTqUWPtpIUXbfNaxtCD9Iebpwr3q7PzFoc7
NphGHFNGoALOAUsTulfRLroJvpYX3bZTAuLcvzSPCeLvkut8QYsBuy9sk+lUZ1vuVumNYc92f6ES
nkyXbNWgznYCku0fS7Hz5JcLyE1yfR9okRT30I3ZFeiHlw7DBFK7L1A+9xOix7OaYbWeaGtgiM41
q4NIQWn5eQ3Evv1WZHQNdsVV9edvlmD7u+Pn9eCBJgLmNpFlURz6cvSp/RkxSeS8t/3urji53t2B
FWsRDnXY0kBrl+JQo93txO7sY123wc6gfNOTIIqFir/A1EkQXo8x0Jssr6qsPXzXWQ6mIDAxZCne
FNbWYKYBVvwkT8fVuWVD7KUHDUH0DPztPNG38ZLqz0FgouWJ/yGd8/2JitUF/awTgL4BPTSJ8Y6a
kmvvTCe+AWJ0rM4XMJZPpmbF2+CQKvfXanMTM6Z/LfE2xSTnC/1tSOnfd840G2VXt3KF97gBSUCl
XU7QrkjDl5hz1gxeAofvTZhgwzdJuHBMzJBRHvtLUyHfbe3be6m+UUrwGhwU9YODTRhJCkO94qfo
1Olbza67lfO4iIdHPj9uj9B4m6IX4cn+v8G92H6WPzaOqYItLctLOlG6EQbMlle3829839GpRHwR
HJzhiOu21aYFNUGfdUHlAySqWa8OaXPii+J9hIcMAgJLcvGMMEOYEIpULNExSZBBg8Q67cIgszEK
8+cbihqjGM+8Mvh2VXUnNCwXk5G0nGY4oHCU9TwHMGkzSeRp/acOtGbfJSgWmw2EAFHFGIV4fKn2
vJqapLXdfU8Y7N0K99iSiBoM6MZ4mfiWUnw1sxnSPsZgLGy8B25GEbt01e5kxdwNFWx80PzTiCzx
pkx8KjZ17S6fWyB+FMwOt7wTwOfZUj+df+YBEJmygoxTcDVi1lfCteR+KKhc7Zov/fah8JsBbY+l
POpTiGrTTsy5YK99q3Huaal4t/zb0QWOnPSoya+xPn0OhaVbvA1QVyPXieE/OPGyZ8Dt+W2HS43N
Uqczz5HIrb1vwXED/d5FDdcTNQt24ZgzWAHn74pxyupknAW7leHJ2aRjDda2a5mvCIvA9vcHyjq3
uZAlqYHt8XLvhPBG/MNjk2FCtNPWxnAv8FWRqcky2ryQFfb1FQL7/3VmwzkWkXOrIH5lxVoRh6ej
6tiMSzqIaZTYqiAt/l1nvH3NWSztoEAkzFFRq83Nap+ef6LwwbodaQ6LHTlcRnl/EMG9Mu8yMci/
/MwI9FZVX7UX3Z1KSwYPYjxgegKEEpI+NPvbZew05kJOcVIO4+cQc8EOiVwcB24Iv96ckOnLFqgr
x9Se2QdPKaMOQhhtuWgOm2M0GhW4ctLBgDVCtjc1PJxhj9s4FBvcnPBdVRZoIfIhUbIuv0IjJPJ4
xkRVF5e29Jh3ElURolpASRqNgUj+wVBCYZ8sQ6ygGVWqDb/ArJizxE5AOJ5a+tKWOvplpAdkTiv1
fa8hfbkJx3BbL5wKWJXT9FOmllzfD/AVUE6k9bPp8ZVzI0GIsC1nd1OwcsAHbcjo+QSLWnMaGTZi
V2IxM/FVL4Jl3aCpiXonOVQdT8m48T6LrxJ/luCC/h2o0T5Fo2HWjCQGfOYggjg5PHagwK29m7FS
wgDUeyw7Z8yqWEIXpuaWF8vG7FPoN7y3DeU9xPzH4m0leTH6tzz+qVZq3AxEUPJJcTRk3U2pg9rv
C0vBTeZRv3C/FD29TJviSB+A+hnjXZBp1rW39d3f4ZKQC4G6d7hjc3RPEozxzLYKNaWJAI5FhTpH
ISi2RtadHrgdbCBWDs9gvztL581cr5S73cIoBywU2JvSZxabPqizFGnYKtsNCSLXf7OThha7Hwrd
k2QpvT/uXCcuuwjn8RArrlt+sGTLZq9XcpodJqoA5ALZnHA2aVFTHJ+ambt5jXcwVMj+K/waJEHn
dYIwfD7TW+ZM08W5OP/gNjhxOWRNSwSC9f446eIc9b0AP66zrGbxi7ypYqiHN4cSM/BGZobvHCVY
zxckhjkXfEfwoqzyg7dbRsrVcsb2LHgtOaqm6zsdikD5op7HHy0pkoqA5aWs7dLKKV6eotjl+52+
dWBlPL5Q8T9ZDRjr7k8EYyFsD1mFpB4lbKNNoNlQIQXA0QOeH0NznEJ09NMy99DoTTCQv7RWCKsZ
tpcE/Hn/dSDaOUPLf22WLyabB1dFR1lkugl3N7EcdRyg7m9LY5s8UN3/QvujUMr/KjG/wo+hSPS3
7PAT4oSNDgDSZTypsdY1w4u5poPeVR3KomVXvNBK2NXQ6cXVWQiynkFFtW8A5+9GKAMLIUmfhwk0
4WX9H1+b9H/eX5WB9P7pRKApEG+shT++p8Mz2QBp+coSxxlYcuLNp5VkruPqNGJEw7x1rGbdNMUL
fwqmhSk+asjUT4rUCt7bpB9aQHtzBnr4B/gdzqGte6cAvomwWjm/1mwBt+Rq4HYut5oYRwR27MM5
GLNqQkffX3n7MYZaz/F2NZn2vcikUCwjNW9rgQwTMIXvHO4sckiuvnvevSlkoYOwOUD194ew6PNv
46BJkdWh1wa+fX1dhV9Pe/J+8CDDZNhUePJnN+2VrcsqSmLHHvSNEuRlFypuNbIvHShCq0vkSb5A
R+RcY7JbhWgnfUsrtr2pzwHilsYjBulwEt6VV6HRdZEEYnmZadAp4wKtbRr8WmJwMwQvY7a7qa8z
mL6kdhlVrIvGhE0bdUTZxZAeKjGZ9rd0aMjB7y9AFvB9D51dDzDz6/it93FaecgnCTXM28z3SJzI
1dZLrRI2rfRV9zf1WcFr1qXreLUt4t2KqjcVVIXs/Y2sKSdsq4E3XZt4kWMd24A98hUQ/f5Jum+I
OYBoYk2dPLm4tto/2N4jNyUECjb0hklnN/TnfEaHPB/VRrQ64Rw93Kv0MxtseC1Tt3jtkVIPyW6N
SQ1bo3DHTUIHPJ0ELhPdwmJU9vpofGI1CpGpUUe9427WabTCOzWi+fJhT2BADkQPTM3Hsy/rCGjl
0Ddsw+7b6tWTAPrTSbXHt+2A5vPbANB/e3e3/E2I8JPIHIjU2ESjfkn0xOnrgSB1hbjQjTqT0cvv
EN0WPXSIx3LPV79XMjpJjfVVqzMHD0KuNdAJebDiLg8AFsiGgcclUyrcb7cwE1C0MgHp3FfeNlcb
wICz3pEbrgqV/sTWXTmjLGYCsoIaHUiPJhSgEYxYwF+Vg7nLoepsVehISd1czdFJtPs+9KRF3mkS
GN8Y+jFl30C9wwanh9V0i2lEvYpXGoADehyMvI4foYh5k3KiA7czPiL4z6R8WYdtYGx8ACJKtOAv
3oK1VB4WhxxLRIPEc90iePekzgz9dHxgjXU40TcZ8jb3dxHWmip41R6oiC/37o1709dqjyXWNM3M
BarJkhY0ZQe0Gtk5bx/vzUZcf0W22msXQWpWExuwmd1errpoXFGX9sSHIodNugD/Fp+s0+eFGP4j
BmRlK5LmcQdtCqR0i/p9+EjV4jSQou+Ht4IHfeMPxcoAz6TjQCPDiScLsNObNv4fVxivr3BMM1GN
VGPxVRjcfcp/ilHHAqaVdq9ozAiQjrGwiYlTpAglMAEZbMLYViSPQ/OjHJIEsasQtdBTyBgaPkLG
tJGidsbwQzNxvykprFeQpVCmJDEtIQ9L+M/h/FRkEhsGvdz9TihA/AlmvWO/AvLLsDf+5inMcik0
wsfGn8cQ2BVyAI3Ccch515WvCDJfcdOGiGTO+0yVtQDg8dT/gSwdSr4A/D6nFcz1/EY1sSCI/jy0
XLihq4KhXYztx98oK2nEOWlG5BqJbMXutOTeHJ/HeqlazHZSVzRFDCf0qZjAt2dug/qbFflExRCC
JFkVz3Nmpg4lH6uVjd80VHIwNlwMJbzZykva2BsCp2UZs+VnizoSD4X3B2qqPmg3tqGf22qw6+jI
YWGO6gpxs8qmvJQSP88UFg9ZP3nNr5UYzkXCve3NIem+UYTGw5xhcQRaWzBpJp6uGYdADW9/XvBH
jdXnzxxHBeE+E6M/OHeQ5V6KEYVArttcANx7aVoG5zSqZdCIe08HUwpZebztiiQV74AfNWcVgAff
HOzErZbxAxoB7a5fBIynSMl0MPuWpbfvAe6C4ppiKZf9EKwFJQPBV6m+G2pT9OUSK7PUheaQn0XA
lSOwMAotqVjtBprL5Q/A/3GQ9i6zZQLRNE3zdr4LYEghDRN8sKAS0f5Bvph1jBuqB6I0SHt5BtZt
eVDcW9rQNWsRe5vDLOlv9m3tzdE4H015urx8dpo+209zy9gB1ueQflNsHrWkoZGK2OJcwRR6x2lu
EVy0XKeLUpOdgrZniIYlECkl+mwKpkC2QgQpARK9OC495ddDh/m2m/VIlpk4EQ+s4R0t7nSxymax
z22HhfHnVQDT9iQ1VqJt7gAci5mqOlrXbZ9QjJ0ww1De3gjUjZvcBPE0o8PX4+f1zi5wl1+8+5/+
DTdvZ00Tpo7/nP3mQFqsazAcfQTyczoY96Vjgvhb6boOD4YEt8O7K9xis0Fij8/Gy836giCCQ8SX
ygayBExmcBLKG1Q659fb0Uwm4meWtK4l5V14RCN5nsQMCa8/4BjCC34OcjnDZ02xvqRZwSEb2eSN
E+PKZG5A875u4A2GQE03KGZwCHetJCF9C0isTW+Zu5viFFPilRrNPLyM0Z+2j9pQ9zX6nVB0D+wi
NODJ1B7XEvp4aU+VTCBZgtrqIfWSRnKbSMRhFU5HSeU7YM0u7VwP+ChwOKIaIFODOWJP3kJrO4mS
tPxRVitfZYD41PczU4REzoaxSnrOK+UM2AIq3YSKNpb0o3bdfjGQthn3CuBXJmTnLro1vJdwhqwU
nFipIDIniTcYjgUHJjocR3LOU+nTs7vuYnpU28qrJ8JHD+qSqIXaqTjqk9GtJCBgtmR5hil3mVI0
EucXAoe2uj2qHqHENpCGd3iLdXFWk9/0GKISOj9g2bWsqmls6argcD8MRH0fBtXxiQgS9dEjO+c+
U0vLjAFFu73hHai9RCECttZ4f58MY884DyBidRCLIY+YuXhSOajus9ZW7JfOdBaSUKBLYxOuOsVQ
iDMWsUt0tP+4gkZeDbNt7yGeweblr+54E5+OQ2BjqPhcCy64Lbh15gHE7/cuEUcSy07UQ/MMBLui
+8zbv1S0lMxDlquh7SoKk7yfVyuPurBSwBR8lbwj+m9KqRz0HI0T1SCEhUgvFT0R++G5Jp92bPfJ
Euzi523qVaGcPkgedZLRTHLeETN2wQXXv2+E2iVeoEDr2i0d9W4g7o992YjvQD7xVFj6RTQxE/fC
BkhWc0sMlwkRnd1bHKJBLSZ2xI908FgcdAZKSNMmlKO25IvU/ydHNLqfGvEVdVvTQ5fIZZXGnZZl
jClX5e/QybNcHQhEiwA8nEn7StOoA5iTsZcs9H81ZyViCIFsnAqeREvYZ90Sn9KFMbwTkQ1oyYYx
ZJCRDt+rwtPKtoUlGp9i8UHAVVt0zb7an30GRsqdljzTeFyi8PVgadqcIFlWCe0zBzmf4JMsAl3O
O+awgW06fhMxbf/I7/HK/WRtqiQB9/Z2AWlEOQs/duGj3YijH+vXixiLcvKQy0gA2LnRel2JuRN0
QWcW5CbN6hsaqaxT0g9jW5rwy8qcQxZ4mUiEAACqbnx1LuUpimFXdHvfYA6SIBBJJUFzkWonHg==
`pragma protect end_protected
