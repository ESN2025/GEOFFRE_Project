// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:25:52 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SmOwc7mg40bV71KBqAhUmAelWGCOzZEWT51NilRocdX97LqdrENoBRhrHALD6qaz
JMr1eNTdX+K1w2DMWTxag+f/Y4r8B6xjsYnhj9bP/gzz28LZnJP9sTnNwaninAwN
XzTblJ+FBtaj2JIo1qnWvQnSCKko2HIV7fT9b8sjI9s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16752)
md2CVGzvYognuXVJG8ZEspBY26RE55LoYCzskl+B0OP/dPLD0VgfxZHA3rsCYWz6
omM+ckkvXvguaYcD7oXltAJAsh9RaZuXikO2eIhLIwaIeBGkWZ7+tQN2AjB0+rF2
nGQkpzVaESkWs6hTV2s0VOxTJBMbcteM7geWHB6vIGe8FjDMZ861XdGTnlCww3Vu
WbeBDrZla6iHXOgoPN43KZgo6esY4QvOOMTgRdCwxotZZo1Z2ucLdNEtsOTaDAgr
EP3c46s8WV1+4Ftft7c3QOBIfh57x2kzGF1qOqXDPGlLF3GGijnwgYBsikKNJbUf
5vxGIoWz355iIdKrjzrCpwIW+zSN4ay8T1I0Nla/cqPcwzB/Yh68rMNjW3k0ku9/
sc86dK5qXeoaS5lxWqMRutZLJTfYM+Z7m1S071i/0X11lJ0fnY77rtNchDkl1pnP
hE/Kd4tGTphC56jF+B1jzyXWmrpvOgDJkiJZcwEJ2ram93W2i7GSk9L2TpjOf0kf
YSsUPj8uSeVQ6LHtxiJA2S9YMHai3PKDaGrwpn7oEN7YcAZuCoZgM/4l0tr0S8pO
kaDQEcDCnZdCivGHAmSd+P3AFYUJnhlOAXFwq4EwsZlpvgtpWUKTSh1lDlrOjhMI
wz+95WRdOnztCapNz7p9+Pgo6GkH5NUm9kEGxMhDNMAwPjPUU0zpmCLxY8AJObsE
d2wK1xnTKOvJt9ZQXiKJ99dw7fGuZU8/8uHmyMNTiveOpmLaKDsv2VyJ6B9lNV/Y
LvUtE+0hCylMJAhkT4Hxfx9tzBs+nWTc7nGuBBOH+5iE1Kdc5OD2B18/LtM4TEb7
+F+YPebKWLxrvr/jYdDDiS1eh/S8Bj5h2SkbEWCCtrv6z+dUSGnqfbPeH6lx7yrE
njEoI3K9WJLKu1ViIEaJo+HQJqSVlBsFWg6pjA1guAstaF9n/OkMSp9pd1jNodle
0S2yvsU/rgWFscK7cpnYASJN7/i1Ye4pFWOrd/vGm2KlW48wubzejFHdNQFNSrQl
3rJmXkAwUNXwEknWV4BeF6MQzdnCCzUatIKw6/WKEwWaviDh3lszQkW1WuHUzKuR
i6DslgzMFXXLlQ5FV69iIYK1jNT+2wFoq2ZyOBQuxhORdScX2C7X/lpXSMi6s7Aw
LoT5c2ZOHppQL2ou92mBPfduqkLwwM1GPK8aEvAUAQdS6ufD1+gFeKjK3GabIprA
CW1ijORphan2C8CKAu1vVdg5XT2tdfj/qU4Oczw/Efanqdxtw9lQYwKD2Ja2TcVb
XsTgt5GeGri2FkIvyTIa7BaFpuFnuADXg2MqUGagz9Q2RrEnwt3H6vtfA14pa4wk
R/MaZntMQdAZPBsk+qSD9FF2GR8R6jr3O103TgLVgOzqgbi+zxkkHf8RUVMwLulQ
OgD8l4kRCWTG/xMVRuCgH3H3a9OHgXJxF3P5Vdw96bqPaz7HtU1dMCsLc0ktz6xo
kJE6T6Mm8kHXYZL14GETilAWRICf3HTegnQUpNX9J/IxAWaguvYY6nXdnskzp8gT
t9OxirbCzgX4eN0A540hZkxJFxZf7UTkJwrInj+SlKHe87hkbZkQ7n2GN2C1YA7x
+bORZBBTWv2WBBBSJfW/j4PDLS0xm+L7TXlz3gzh6VbcinRikzlQgyYYBNaNSgXs
raZJqjyCt+GOlqLm0sF96ClSjRodXP6Vu/N16xIUcYjeS5IUcSR+YC4OtZrEo8Gw
AnOGhTJN/T5lJpL9V87QHGlNOiWqR5i2JI3iORYaDXsH8DkcLxs5F134uDWFjNC6
Sd852nANgAygE5jgrHqzrNymB7EN+O1fCANwcZPAJIDZrwY2biSdf67M/WWaI8Va
YIdCglJBbDpltuTmZccgL9YYGvEFo79UxWllO62J37nUFFdSzzthtW8r+4qOBzNu
8vuu023FtRxi/1zHsZJTZhj0vJ7iMCjWiW9Cwk+WKtqOkvMz420FMvMl0qrcTP9H
3K/a4lSog0AcdKvC3z77cytXH4fwf69KcXV4r1NIrD8W02FXnJ5dL6TSmL3mvyLS
eKj6+SPZJ13hHGi7uC/Tgf6K63Em+6Ur9sd9E41L2Yr1pkBWnCURcfP5/BrDlx+2
AhKOz8pJem+xqkoBM0Yf4wRCSMY55FvnMCCXAsM8KaWQjMa6SjzgJ86AulKfF73V
T0Tpxkko7xFxvOTSsEheSErmabukplUbQb03dkmeKawxu7GfuJE+XKGJneSy0OlG
T+o03+CO3i6KY7saNCHtLtvdPw9Q3v4VXbgHQ+ZPL9zh7vSI2uN9cx0L/g6SJ3Uv
u3O6kFn8wwRpQkRuyhJp5LxC6zNJ4joA+uZYTwiysFk5TjAmKANDKP6UUWxNAsTY
68jTqjDQGUMlnJYhXULpNNlQyzrtmeqWLYTMDmDKq1+ejSpfVuxfJk6QYSZIbSUl
epkh0MowGCUVQfYjjhqGDboxY4T4PCkdO4OmmrgHIehJa7Qr6nVyNuzYIsZDNM7a
g2GmhcGk+PK7VMF7tfRKFuIWEDLHnegwdswVfY8axjugnZ1LVWzdA0T8E9t3ACaC
3zmtHSHS9JbcQJ7XB6xSo4OyCJcd6JeGmg/UWEDSRpTTpZiDYHkHufc7Za7lPHQ8
+YIdTzMljrVvtgzjxE8bF4VhceB9rNutl2hOXUVgpthAzbgVSM4Y3zo5XPKOlWcL
yHTHur+pwLqkWMtkahRf6kdnnPF3qWhL5TFrjwByFYzs3tW+iNDAJ4nkhZK8rTuS
0Wb0Q8CXJIyJkktlTCgooQ9rwBLtHWjHOxIJvHDts3ub29abBC6dx1aVDoEa3Xuw
UtIVIz4SCVJLN0ce3ybmtdiVrhnoAE3lk/1NKECXGJSoUa1jh/m8DJVy4kSl20VZ
wpVGKk/ihl6UDIe3mJkjsV0WUCJvp5oqUjchrJFYkMZlds6Cu8Tss67fvgZ+/PwT
TueNCXgfNEoSUCZan0GEvCBb2rM8FsoATx3R1cvpLjdFTJ1fBzBGiBMoi0PFzgMd
keqm6YqMd87wqMomX40rjD9VHhNncDrbGvDwvkwtazm9Hlzj/qCfqs7L1++EIVBt
gf937vCfqKyXOk0MrfNlZKSGyzkNqTrQCAwwBLTqhTQyeHwLfGa1bbZ+Daf3KnEz
RmoLY+tsC9fvMDf2rUGewQw5zb6B3BNqRXR7BbBpoL3IlVb5FMW6xwgs8ClrJStc
b/LFlWx1i6OQnNBOx7QTAM8QbIKkG5B4r34YW9jngzn52YfMNo8fqnanmTqX5wMc
QGmPTfHov8II6i9nr4tBhEGRcTGoHmaOoS1BXoGUGht5zKHVaZ1o2COixbRB2ytq
OWE5XO+Otq8moiHqnYYxFbEYuBQVaDF7No8AxAkdR4bhjBaaybhjoxaM9e7I4go3
vC/yGbkz5Lyho9N0V5u++7ARBItndUsQxmwsGLrKKn/5+xwNrcdv1EBG/p7sNMjK
U7qE9LVhxja4K+UMhKxuzGqZEmXXl/o7HqmHYRg16wDnWHLqDgCqTU4nmwRZg/jp
dKeIP3MSg03CdcneosV22NNJQmc6RAJ+lGBeKiYmLVkCQVmPtdoxGoRX2gobR6zH
XsWlCZ7K+gZ51BO1nFLHCC+ON1w5BEHFl3HDFqIvRnm8HIBM8n/LTQm/BgKjc9xD
ToVo26iy/RWaOIsWLW87dBIjzw8wVKWwztK/1PCE1ep75u+gM/B1UnrzkF5Rl3Tl
4mAzWoEiL3iUh9K+jiip/NUkRKoxinQjWrILiU6KBJakEaNqRnBwxcgmSdTcFgg9
61WfeIl02/LC9rsVdB30W6B6+eW+RFNui8A63I7X2KOHqWYM6pUcv3ip1ztBttg0
xzbpwowJKiwqmzagIxdy937KGi+iFCJ9OYP5JUZfolq/H1SOcw3iPyOuKxt8gFSU
VgMgyBdYpVuLXnwhotK7Eckxz21gpdWZbE3et17iR8hJUfp1/OsKZ/C7w+E/DZpk
xfowVGDFpVaHYSow0H+Appqrx47d5qllvTY8AoH7px8GNZ1G1tUOtJ3KM8BQiSEh
qWmSZtfgNa+0HN8GbrjABn3KAo4I40zXCd95NYeNcsx46VFOnzCGT72vFjLMt1iL
nK+Dsb1uu6FENsUKm262nYElzyFXywTpFkxlvz1BUI64EBx1eG8uo+YvLFP2uwfk
ApxpvpUZqsmx2y/0JciK8Qc9Nv1q51DJzrgbh7pyjS6KSlD40n7fkmSKDgRavYYB
4d4LERfxdyGQHlYzoVtem00BUuhDfYxCYebwRpP4p5ZUwijiuGv8Ry0qtkfUxgN1
6vBKyB3KjzgVGc8QNPaftg/qqNwxIzJoPPhsA4H3ZztB9RNGKLjrqJCgIc13xaKx
7yO/EjIk77y1Ha89TKnN4JtpMXRxkldYpQ9QklEaMbVONGknVjjggAXjTO9SCNRP
2aQ5q8Y1i5z8TF6MNX7Ck6QX018aowQZbJrCC/NIdjtc+doNbJ2kthVashgYfj9q
6sGlFymLxhKCH9D59qtKaVu5yPO3/4ZJBU10yvBxHJ+0yaNFbp5ES02NtUe4jXwj
7s6ZArQMtFZZubfR3M0BEmDXzQS6f2XZ0wpMu3PuXCDWXuRusiGLZPu1WDHHsopU
6VFFIMrwpEqbkYFzjjLa/oSbXvFpkdgSTPQ5skdRLnzcFdzQHENrRVv64XGBEFTF
GVyQ0fzOmaDAkeUcv0T8WAp9IHu6xLpbXn0yOOXOSHcf9t/B7JrN7ImooMzCkYOe
dYUCAmAx/Cpk+hVvZi1qVRoRAXtH+jLXVWguJy0MghopaKbqvZz5QTLNt5Tah9L+
zdpjELwch6s/lgT5VAc5+4i1zOEbiFrLhevFRnn4A/tZREtGo/mz2mHGdzQ6ZfJt
V4pHsTJzr5LaM+n/zbD4IjCrB4NEdGWwE8THjrRoEe+pzIADNRcx+ri8V+O79Uff
Kyvm2GVjVSVlbMXsgCqDJ6ggq+71Xhc3wTUp4VqcOneLD5L/jpXSAm7SOL24XIEo
HOgfV1yREVwOzhg7AzMGydvPV1JiQwrPozTeFrBjJDf/j2e/dAXXL5qvNrNAA6u4
jQPVZoBd37NIiwlQprs2zVjug9RAZZjDJwmjJUBt+X6nF71T8n2BUbOrUT2ykHg7
/6luXuUDTeAyH0Vj9CShJlVb6R0TkqRMjZKChUkm2JU9ZAOPEJtJO41HSgap0uSZ
bLCjKrP4QPknF0NAd/+bQi9tLpBgXOYpQSRI8+dGjYEINoR25ZY/3eklpvI3Qbey
WUUA141jJj7D8DBelYaHN4sntOUOUe8xy6Dz1JdB8nRQFjO4auyudCvSUDl2Ar70
s0h7dn60SgTFNUZnjRvJ2Mn0wosV653caT0C98OaQ1Wgd0S4O2K268yq1jdvGp2M
yrf8Wx30BixFLAHgR4YmL+TVCYYVw593epknhhFHyjldSF9nVFPdOicxmxGn8+9v
/cKQ3YIjmeezoJz5KjUreZ4pxLFbmLn8Sdl/QvO/3/n9XQTYspG7ApMTGPedG6ub
1dHCXg1qeJ+BZvlp2LSQxVY+tNz3QQ068S1+KmLH5yNoo/l1C59JE2dwNXQuoDPq
z9pR0pJke3uQfYuH5L4Jgwtqrpuz0zn+5lWbVmL/DkEquTmtKP4LErvZmVB4E6Py
D90MWC4do2FGRLoFFH+MyJMF22VlkFwHlqw3C+Oe7dw5qrEEthtyWYhhvzaomfEL
omZOyhrin900+KnoQ5lYFPuc45ABxgfDpqR1WUHvYcOUknMc0HVCWOs2anXwOPGM
CrZxTAiDrMj4rFG1plkxuIltQJ6P93qyfXV2kAm9vcY777FTVRH5X2yx1epAbhMI
mBqPat+44CmlnaIXfcEAQHT9UQnL55F5SCVzYSf68b3l2tKmUtEJbMkPn2B9vpzK
lVb6yojh3YFS7t4uPmAAQGv3SnJT6LfByeKmy4ZToawe/WNKIX9/TEysDXBZ8+Jn
f1mNnxOD21JXElMy6sRuQtTAAIisAtKWNplZDjW4Qq2MypPUcgQ1RFgAsKD5Q0Pz
51MomujB4r6T2M14x1144ZoBRoPBCkBnKeTuszuwtuJs71uNtNEZfBqQjVw0DyU1
duqbOsp8PB+Ub3Vf8MZKPju3D3lF1TBOqmEpH2cuSOGU7fbD1b+OCg24ndcTb33E
KAyO8R93wPLUmdkoT3e0uWrML3QlO/4tTwd2VcfVVtIGyt05i6Pq6toStCSDcbpI
AmrR2dQB9PZs4j7ia9oHSvjJqRk0a7r4QJ4/wQIhzSN52hoQ99jzCTFbkPnwEGup
dY6yf4Obt+B62LeRVVwDvGyJxHTVG2maJ/v5vybAWJqIzhTvFwwc/OxuB0JMGgzv
GT2guEexqX7XxuGnVckJge75B+9D/y04dD7jwDZGvbOP/b9rUI3G2K7ZMwK69Y8E
sepxgFNZmC9v371XFqQRCZgDw+srUv79BhVOP5eLKGec8PZZQH+HeNPa69ECbQ4G
6R+oietxAdn+ttZABnVBM4QM7nM+F7Q8gB3wu7LGOuEUb2Lz6KwSzdKTNT6Ux6a+
Mr49NTMpb40CvJi/lmxLRp/qpc7rCZQRoAtmhbURcNsQ6R7txFkUjdicme6sp/fM
rNUU1Wk3nSTvCzDotjnpDIS4Fq+e1dKTtqImNvfe8sSBubjcI/NWN0gJ7KRF8CDU
+VI+q0pMxnr1VirU23vpurThwzgSmhBvdcUIEVzZeq6G7Yp2F7eY4TZASW5arHYL
UPlgFQlHCoLx7nRIGIq+rajtWU0Rmjw5JkUWGnYrJp8IW7qjYd12+JaOJZq4zf3r
xnOyF9iAQYtfb52aRxpZW6nFbpchglaa8AeED+e4GsRwcPJ+LkVeUlrdLk1qqx8Q
Jw84UDRMDkthR6CED1ZBTMzbi2/o/Jq+7agaznGaIisTZK5y/VxvQqd9SiWaA9aH
6oZo6nY9C/avrwHLsLqeLifmwW0MyCfC3RX3nt1FqcnPAKzwbIhYE1tnmQhEAvuP
gjjEZMP0lU5M9kRu0cdngXIoqqZN762zvlm1QPF40tU9PQKj0oa0fQStd/nmGVqt
9GKsieaNJCXa88DoQo9SS8jKb+By13SaBKjeVC7h54blWZC76Uz5fBPZpuIKoKvC
vjjYt3K9B+d6quOXfdaz/2CfHA0Xma+WNtSpgJoY0FHRjWQjJoNqAC4gqQh+0/zb
hnRwkHyX9qQ3FUkbHmxwQvqrnj251bNO6Ei9A/WJPm4YSMZUTCpcQcJ+HxGWhlt2
9gSdmUVyUcw9mv326KTe0ibkqNOADmCNb2oZ4vN3VmS+vEZ6qfq34LpADQCcMUE3
Hx1mlF4faarm/NCU6x736VBaMHuMWaB8IHD8KHJq+cwC1qjZRA7RHyvV+nuRZx5m
T2cCN3wTiAUTky6yZh+GLZQNSgTsrq8yYGx0R6tdAyV5iW46rE/4M3dIVPPIBQmO
W+pc5wEg3ftZlL6cO7R+cA3QbRsE2JKu5KA+aV1L3+AMU5slkxFJ0d6Hmp35aZn2
mblF9O7T0hBOQ7fulO+aGJfiullBTodLcfn51Ul+C8VIxIbHZRyEIVxGAwz1IG4c
DAWkn/TybytgsIyc+nmWMQVjt9Tg+ZQb3U/ePHPadkHMThR/mT1ypygpf/u2pPqx
JvKq5J7faDfczZreKisfdOgA7uvp5h39n1ooVR8r142ZFT4Ulp517xrviZIG8/Dq
X78b6e9V1dj/kRUoBNVAP8B8Sg7OzEt0x/rlvvr8DlsOlSrWJYsFoxazDmxP2hHG
48zwi91QCOY+Ac4TTyAcX+Gro3UBaH1lEj93HJqJxwjSDbQd+N9qgQT1XucspU7G
Gh2x2KB/di+9xV16COTU5+0NJ/2NF77sMMybLiYW/ot+062z2SKXasMqvP8mqrdh
2y+Vq1+l7aLvH/pBbCsvq3rET0F8KjaF76P1IuksUiBeK3a+nJRE5ebgHZb1zZJQ
jzLL6DW4/WTxZrB3G0yhJfwQOtAZde1eGe8EjmjERx09/Fgg0uExLHefnWTzSeJA
RcilM5UeeVrQzAIeQl//b8FiibPjRtJ9Iuz5cB24DBhXy/e3pcvw5xSNIAQjoO3w
vCXFdv1ztZWek16ICbQpkdZQdkGIPXnYEQMof6le4aMHrey2fpC0tOuxI+c/+uD8
XeWNDFneIsDox53mMO+rmgSLwdgmN4rEp/ilxGMu/Sgl04xD51R0ozNTbqze4LpP
9oOm3m5Mrw/aibzxbRuo+gLt/5BmusxPtPmGRX8VUJdPE5NYBwJIq7qvGtKNW9NF
m25lyNwHbJ4C2ulhqCblMXexpPi5Ync9NcP3WJY8hNq+q1qnJUUTc2SvFUek8w7p
Y06+CZ3QEbRo0Pf3FArL7NTD8E33XAx1VuNZRRUq2c6cyE9Q7EzRNKPr18rbzrYK
fevq8c5Ht5Dq0WbZOdvZ7U122j52QfMwrRfqt+lkxeFus2NVbVYk1YC4clcnoTw7
a3CGCRyq73jAtxkK5T7RNMewGuXw1exszncJ2gGj0kWwBBG+oqF8oLTR7VopY/O0
HyG6g6SzEkzhRxj8osS3/QUDj2//+ZFCm6ejc91uSinYWS2B/2kRfMzWQmmlJQ+9
/fZgbIMkdI0d6G3dgaUnyiom6Om/QQMckKrtXiVe3qniVR2SqFzoUheHq165i9fO
WFmn+b+T7Wf1EPgD5UIfNZnH9N145KMGdvj4HLi69+Z/6CtwU01kYX2l+PlqV/ke
ffDCsROLoSK5fih7dAAEr5uoVF1yWMCn5+qwXjZ6HbvTIVCbqZr0an6aDUCW/Bc4
LKV4ndJnvAfwPr2qaxsU6OASlWN1ic4rwLhArg8FsCu5OFtgPJGTcm4dnjPNcg9a
NZW02E0g8zqmSvSw3N6ei9rcU9TGJW2ESdEzZHjXAqW50at30R90Fw+0v04k089l
FDzPWEmqnNd1Fy0Ar7wf4ed1HAPTj8vpmeD8tvI0K2I1W2s/P8assIvPwsftBiEI
YPiIPeiFbW0AV35OqhcMqRKOHN6kIDhVZQsakVs6LeInfso20k9/YTeahhfgEd5H
moSO7Xsr11GfAhyywZ2Q+qWS8rGm/0VCwrpu3qb2923AdDYhvbSLjm6/5WawVKoZ
rsRuJLB/QjwtMSIkP+IF8tLS+MGqBYvoe1B5zSxJ66oQ9P4exE6tp72q2/GlzNrG
CBtLYbqfFctOHHaf1c7xZBMt+IDNnSWnsQLehWvaBCTElUq8HZygSq3c5CFo6mv1
gTw6Og/WbkoRwydbpK5i6nR8/EDGFsguN6cuBmBLoqKUZttUtmNXaK79ZrtW1d1c
qHSkjOnMP8Emx59Ipojhv7G2VxJ53V4VAug1G+MzbjTw5UsQ7bExFgcXGhDFhkxh
9fJ5leU8nirZio5P9P7a1MKPYY8wPcSIYIZ0wPhhE15OeRsFJs7J6iOpJicXuO0s
zSlJ34XsdVmW2W5p7ZLbn4LZNm6rKDVwzH/zoezWT6tGtDNM8WP4JRsHiXqQzim6
Ny4zf//wDhtQlzdHe5VQNxevO88laKh5qPeIoPIEke+Uduln9rwCARnF1CYaseRg
lxRo2UMvioi6EuwPMnQ6LSqeLYjfnicD/eOfBDLDmmuxVz4CfJpQfc0crbE4JOIN
eOfzu5cOdife70/oIzXEIaVIziX/TyoQ2/clhCpF3wwq0gIzOBBf1GyLiB1Yml/D
yeSySgSPliBjbAVl18mwg/TgN1hYxcSxHcys5hWeXY5d0RLz/FsRXtW/Gne05Krj
rKAmVWI7oo1u0BHde92tTiENsGy7Jfsc8Wc4QNYnNZPdiEd4309NG4LcI36L8Lr5
AmB3rc+XJoz40xozJFDeFku3NpNZuZwKE4MctD99xzsQhZL5cWURkQToJLESXaxk
2b3nBVKyikLJEN5RZaxbKUTviqwl2XzDsj+eJGeXniGwM1i81QMHdnMTHEUrnIge
8u1HOL8FgOWRxizIG02iDz6eUwvHpzQs2H+xChlc4sbWQeJOphtxmFsEclsfyXWw
EUyZWOOc5X6j24LWcnS3WvgBQh+VJHQH7PlZWpFY6m1JBtW+W5LCAW3IPY8SU0wU
FOPQWuUWRWVfgF4ElqkMF0Z6kKm9cOiRHeQYJDZBxDGJ/McXolfG9vuV/2vUi4Oc
/LxucMeW1Xj/bApXzyiqKt7TaI/FC3N2pyDM2TQOuHOIvu8aneYScTDhJ8yVzO+0
UwHEGYIWbO6FDSfRQt4i0fnYRPqqsgw3YAwSfGSSaLzjZVmfpRXAslMcSUd6mYS8
46kNg+t8/puYHnRaWThqmmXFOlS97rlXbv8HtabZqeS+HGya96g6/7JQ5Lg63Rkk
OO3oJLDx1fL/ymmOFw2THf3STvwbNyaYzsVlz+6vbgrUqG8+T/NmsINR5cZR87ia
s/wy9EwQ1cXMMR5prsBJ0ZJZMS/DijdEYKXcKZbXUzLBpWFsrsmb/L896msGWGNr
K0b/lebjjNOKTPaP3yn5IAqt0X2bf1skp9AayM2bLDJsGjw1OJzw21Iz5f+sYjKT
jQYxhFrunES3+fJ6XnCoI92tRmgHKZ4bUDhnlBj/uZ4Y7QxdcsREWV+a8uzztaxB
+cQfxgClHQY+NhbiqE3tWahe3EtuWFUzgQxD3zAfZCd9tV5Mav9m01oG2ewZgiGp
sk8brD4SDsq+qDkuWkcgZjrf1O4xruyTqCGhfnGang/pf/CYZRtkR8l2I6lYbm0b
2u5WIAC0D4qwmvazYdhLtdvtv3i31ojRFwxcE6oRa+6G2NaM6qDN/dUwCZujj7MN
cUEKqVAXi7Amc0Zv0IGGUlBxGLjL5JitaR77cXcm0vz/c5Qm7poJ5DjEBAHLdLHi
axM+B+thVfIR8reNEatZOXYwPR3NkzdkN2k7WQL3grUrSPuxMbxwnNKfwZdHLi5n
jtaI6Lx3NFjXWCEnrgRShnUYS8/1J7AF7jrQeD4mkEJrgmqFZGrRlba3gPjWDH/p
wFX6fkNHnlvPr9gcdlmbGMeUu3D8p188DWhJEphdv8+XK/JS51GCrypJ2FxeE4Il
damwGDDznB3l5aPp4+YaqGVypwZNVrro8DjJc5/GcsCbkfU7JYvZfFE4i04F9M0c
09hYrNRPuNdmu8gQkpPtXw+B6FfPCF+ibhuVLBGFCI3WAMrz348CH08ts88ZM1SH
dskWY2Xi2lLu+S9Ja4V4Y1SpVGZXVXuMGSU8GnO8blsQ/rgYM5oS3HTQCRcgkG3L
ZfvxFivmoo4rqmp9lO17r0KOq121Gk1UOX8e91UkjgDitnTwsAWmbDit5yeOmiV7
L7Zbl0BAsEWjaO2L6yLPsTxvGPprmuLl7uvg/LiFj8ATJdNU7J5gZjnxOOq33qGQ
b0aOJLf9P+FfNm0jQ+MycyL9hfb9eZysdcS4BnqliQS2FBBFEbQlCF5qWs6iTrMp
3LevM01xqj2Ui6WoUePeDyH99qoXWq2mBNOXjrT69eXYNZAMMA8MmZnhhvH6xY9J
T3XG69F9V71k760Q8Y1Av2OyJ5+Ql2dZnIYhEgU/pEZiA3S126MC+i9eCsy5wJpZ
08b4NQYFQg+Ft1ECdSMXEJCVTG31NlCTic1x0OBM1SJOBooipnAGMs0lXZLONK4J
IGVZ1iNLhJvioNMfQFzKFW5wRIuFn8veq/gW/mBZxQI1LCiYt+Xs8Cl1yqgac0Bs
dPPf/El2QS06tjPYHmZIDeVYHWkzwHHJAfQpnI+11DoVZUeZFe54+3S/gGNT+/mN
4aYGrpevV93S5rJ1penDd18PoVU4ciyBiiLM6SW9iBj09lRVywvLB10NzkQwNQFW
mGrsi2hDVkbwSt55xampPFFdIYpbbt+zxfAuLsNAp7ujvbN4hL1/Zp8Om9XbKcOk
JibY05dI/McV+SDfG3UIkmFf0ic9lVco7icB09Hqk2MaNHlwOzGORag8lDh3r+0D
Tr+H6e1gzYCUmeIyvQbOwFbLrS2SRW3qXnt7G+nv/A3eR7iJJnVZeJBHR7Wg+E2j
ycRAFPa88tw4NpEKcOdVIncGIyG1fGUMACxCR8QDdLTLcDKq9XicibkfoKp33i5L
2wMUvRLMcmxrHuK6H/iprvlGCEne3g5Abwp/6aL0Jrjwzw/ACLYSLEVmpD0tE4KP
CBvDxd/l7SLfHuYgDCVstdrkmPvNawZpp71lEATuGBjiBMKwPwWEmsbwyYiO65gN
GDJmUMJdDrfWIilWQq2mfWaIrNnzzjrKanxfOMp1fKBGMxXphDZ3O0ZlCtzAphbc
hs+tvZUPBufaRQYpgEq/wu84vNn6woYjLlZ2oMKQ/CQWellmjUEwr8Vn/NzQyNNL
EK3urJEUge5RqZAgMXRLeStOw7CtxxpSCdveEcWX1Wtzdtnj/CsX1SiSQE1lu7rz
NdJAGtIlUYoOHbIXKFl3aA0T/aCkJzRWd7KOn0PLJhKTFm9pZiei2kAPAhCBWQpW
1NcPXsLzaNQKLh0ECvZJOIc75owEHAeAi6bLxmNQkE2BwdyICCS7RmeBj+obf9Vl
29s7Csmc+XSZY8kZpU3TVftSGwaZ47dgxxfrOmB94W9+ZEQhHYK0hvDTM7K3Dhs5
ju8yQR0dge18jftC5Xcd57k+47eFG1KAqjGbX/5GewoKt6LSVUst9WhnWXMWP6SA
1L/MOHq+skMp5gqV2XaP2fxqO60JQTc88WA1ecMAqp71oLSk7G7R9n4DCNKhQygW
M62wJ+/X/BQ/KTymtoagu9st/vrry/VBuEdCq/GLDnUV5LjS3WC87e6o6XTmX1Qp
uRO3IpcKxT+D3IXoGOn8208c4bQKeBO72cW0qOf5KT8ozrKQbMI7Rab7bOdVNiPh
uAtJSrVwcevpV0jYED6F4ptHofoED0RISL9pzpCZaNg0uQcVsL+5mfOwR8I32N9F
Svl9rj5J0crQ5pUhUidISu4K3twtsbLqQyKtC2zl6V+8LoFCbKEG78Iqb2hXZAzG
maRF/Gu5ErPMnt1zy5uN5NWwQ8Ddsct0bIjc3qYK2h/byqu1CG1B6va4WTqRyVVH
NgkhHUK5Ti1p0+OQdMemAP0j5CkKgLjGUwcIggLO/JvoGTi+Z9iwI4axknJRzuHn
88j8faSOyUjSoJlBiK+r0MnuxeWEwNWWWIklDGhMIO3m7W41eD7X3CeYOjYy/zd+
lGIKW2LyEnMg02wgAhCmnq+bMI+Wtg2CcVLEGnIRaD75hRgxHukqF5YZJDz6yI8y
6zUHUa9xO01i97dHbEAPIKMUIDodFXY+95AN+H32O4hMJ2y1Hya8KZeuHX0OGkDr
Oq/rzog7E7d8g4BNXD0Tv+6/BFOdb5RM8duSBuF/x34YP0r4vme/X+uLf2sdWSK1
qLG8FLAJB8TA5kuj+o95YqIIKNwpHXNLFGbSId20n1nST2KaPgFDuNfnS1QOoMr9
hChx3mV/nKzoxT5XPmxFc7Z8RPa7/W/IxZC6cFY+M+NnefPWilWLkJJocDZp/u8v
iC9f/wMwtbOm+3vw88Mnv6qyMimIkHT5vyTlHKbQUsJRIHPUJYM5x/+pOqm9Bj13
IlzEjRIlZ/03Z6by5r3h6GUsS2Fqo/h4gAKKaxKBMAmG7SDOeNNn3AsPtZ0Z2EU8
PkbUZuS+3aEAPLlsLetHOC6qoa2hUtOlVX0DcrdR5AwnW1yUGSLI/kDJ3FfKWp20
Y9HX+LIlE4rKpA4lw1d/3RMbY1RF8ClGRWLrhDgJRMMkKxy7492PB18rUN8pPeXx
B1vrNL/pQ6aMj2457Wyoh4A5BB5K4ajKu+bP29IifPQwfZSk7js1ZtgxSIuEe/jd
YJ5IvpxT3PBEMpKxoX429pcf2b+ap8AkWWuRhuckkfLfLcs8oLQqY7wcBQwsSxTf
UcLirJ82fAszR8J86IiklibnIwb7Pc/9jeSqkhm0g0ZEHv3FYC8wqSVCYsPBoeJU
hyH3YqyyW6Nr3hoKS+hHR1zaJUe2oy1G63RIHJ+ZlpACLQdIe8Lh5JPz50oUweif
6vJ7ikO3W6VQdPZn744KdyDXjhAtIGer1LAdfzP1u8EBdFXCmobgJgwrLWiNQ18t
E4GWGT7tB9rsidOvkpkS3z9IzpAoMDoCaKRZ+pnsTFPtWCHpPxqrb5tBpQdQILTf
V0H/D6u4sc7ExOe5MvrKqgACgRycBM2W17jn0dc4Z9x9+pA1r4q9muWKU1T+6Z1l
cCJPS09gf7JmS0igFhtZJCiyo0ouRuBOtOOCtYFQfW67xU1uUy9Ef415N/VkJhbY
szsn9KdNEJZcC29i5UofWvtA+qypsExDOUjmjaDwZdU39oSFlKNq5cB8KdwXWGu3
4ZCPGOOai0rsDMiYzdZIX/jyqYOMlSEgSX0r/V8UjSyZjqP5LBlX8L5exhE9ospw
c2mivlM6+HKVb9yo98vPYu/CCi2KlRwMWXA3LRje4U2VWXaRoil4PAEb6mMRImhV
JJdtJzFJ7XkKJmZp18kBqcnMNvkngtcXXjF+AmN/WeZuPZ5i3mk3hpcyxcTH+BAB
qCeAKPepFUMYojxCnVGIMJDO794K32f9euYkzj/mbgHWlPoiBf2VlVVZyyleiyrw
DXN3L0fwtuf8kXeSSAoLP8hVERcdQl8r7Dl5gTbhPWLnrTiGwdXwEYxLH5IoZrAz
JrjLsyWewm1D9afxjEVR+PoIqbWWZLDwYadst4hrM2tELkqxthiVbmzvLgOiYsXe
fhw7sQnixK5UCXMIr+I9/U9XGgOazuyIbGttughAZ+dqmXCpewcT+Vat3lMTKDwU
E2P2p7wlB03TXo4yAh4iP/Ki8pRwiTfZz+toTNPaEFOYNPBqY7eRciGiCpW0f64D
evE5mActoLUGZHWA2eOqePa36rbUpEYDRe1hQB7/RX6XOwfKGw0Z5cNIVLIXnqFB
BGdHb0gZ6xcTg8uUaX7RvHvDwRkEdJ9W8g3S836AEhQKKaCmNmK9jRS8HGRVxg3U
2sWrkNUfUZ2ueTjhiGzjGqqae7YEKVbTvSdrFEtMAX6tcnQSmC3kx4MYVcbjlO6D
XGh/7cpfgvlAIXxv+ifO8K1kLALdbvwX1anb6rJtEE343yxlMZ6egNQYwDsiHxPY
uvjB5kw5lPohi4sZUAMQaeT1JoE4oGvPXKfoAQ0xQP1GkpQ+JPbaxyTOCie1DDnW
55RNR8SnIr2LTidPHCf8A0VKWifNdfbM02/rwlzgySp2vec4QzCMc+XjVfYb58O5
c3AsVcGX0U3pCLkssM4hdM51nqVA+B6MQZi/DHOn0Jw3m+m9XTTRxrkNKaH+dCnu
DXvXew6IgMAGDB9dxhct5q5AwXG3Tcpy7Oo5YlsQVvZVSyPqe42YyIC2fCSTE1Tv
fXQw8f/KIha6pon1UwhnP7Zj6KId/JK+K+gdICzDMBwAo9Q1UPwQwPCE69IRy0Ow
KiyeQgMzTaRAt1k+7PoDkrgoRCcH+E+kWTxd2IZq7xGZS6uYoE2RIJhAtX42aVWh
CZ6XwWKM08WcSKgPCvMD+s0qUgySzhVn2eJ+5P4c3N/Xr3ZckK9dfDeV0XBNjHhv
pl25Js+NViqaoyTR0lY57PgzRRqj+lMpkYOnb6DaaOVMjzzyoUPITvM/YqaxSCuo
XQ8lly+yuOohMjKt0nJdsN6y/drwJ6dg8d11P39iIFg0HtoflZYqVh56K8B2kIlu
VqedvWoOE2WCtLgeTqefglIdXsjbgGPZ2e3hO66QGYrE4H1+J9m3F2Oiv119LYQM
rn9NkqEoHJ4ODaBvBqf+hSGAWV1yNMy2ahKGSnVoG3HkKf0E9ndPgBtQ4JRKJz/t
to7hca0zgt4qI3uLfxhLWKkwVsVxVu+CzefwCIA0U9tU+xfxFJhLMwpowelqd2Mb
sWfQO1L6Of93ZhI8swdXuHM5Lei9NynQq1Fq1dSdT2i3YcIGv2z5u0b5DowaMQzb
N4U4kpT+dKCsyeNeX3Z1CRy5vxSGBIzxxLea+WqIpqZ575K/g3UdQkYZRPzP1Oje
hHN0RhZHglkm0YrS2OFOybszxhnQE1w34c47JnuSZ66egKlxmDxhLAAxEuRfOtVj
nhTNxtMlmTRmGT5EKnTd3sXazFrfGQwUpLns56jmWDx9GtyzVAxzS1yQtKe7V0OY
lo/7RP/x2uJ7SyJd4V+QN01/NC/QpaEJp/qOHWl1A0UKCHfDpWcYJA8to+Ss5RLi
AcFbF6Jnv5xn+q/8QM7BjpUKv7Bfj8dVoTk3I3Q6DAzJdMFhj/MXzUQ5ukesrdfQ
ZzhcyCQkBc0CBLK6jkmcKoVFu/8rrgqvpCA03nHxtrqplAE3aiNNhCYxZdwzjqwc
LUel3Fd+lV0+M428cHrEFiftnAW9nikMbk7X54SQg7TvjUfBGGIEpwZaZ5QbLagk
r49jReZcHEeMEFXanC1gyLhMqItTsQ+a6FF5HCiA7bXx7+SRZnNL2u+8r8+4l1kr
kYTbnIEVOvyUtB3hWlxM4whHiuX3CQhXC9M5Evy38j5bJdT8VllD/x/3vh6NfFb3
2IPbxgdDOUmQrOZCYGuClMT/5h/PSyRiMYfGYfKwrhhL88gRHDXNnCTOoT7bv6Jm
4AJZuWWAmTb+plzlXJapFHeoX/DI1aOvOF0iMvC+UlZSxBLhKcB9WxcH/U4ZDwJP
AIH8L/78UAwhR86pZaIZbQ3sF3KA3kgL28uY6Kn7M1w7XJRX85X+IUZHBaLrGCjw
zKnPjJd/Y73J/YqiH5Y60oDk8VIbjqkzR5yd698YBCraFydQ9aP4RoCPB0/l/CE3
xhkidZ2XW9XFKfuuMGW+ggiGoXAgjo2PUEx1ST3yld1PfwsIMhFvswKaGcjy6E80
LSpYS+dgaSoW0gd++E0krXXBPhYSQ4+gsRqrF5y7TTHFnvZA9Zfhvdj8Zr3oHskV
GGjeK5N/aqIppTnPdfXubgpT71wwahEZy0NPlg8kVAlRJRpbsz1mnX85QmIgy/qF
RUIdVBiUu2/qqLlcPRETGUw3cWupn5GBb+BPCwjtkxyQ1/tQo5ZcOtYAwLqmbBRi
6+gOP4853oNZXUtnszwXNzMXKa/qU95FZmCvqwTtAGexnSIvo0pNMMufv4KvUrte
X7jBUm7C0gacLfrq/gGf4dqMuFKDWPXYq2t0EvKnsLyTo3K8iDvhJpms/Wc4iHcV
5M00TPqgjnA3lnJYnR/QXw7JFjiLRLCs9xBJWVJwgLXTcYSazGmjgDmgyl6RTs3l
vc5gaWzDt5QpH1CY0EuC/i/3id9SzRBel3cwwaev8lotmhfFpo5dwhwEbpL+RFE9
zilI/Lv1tDHEgp1+Drl1H7Y+wGF4d8xHB+kMjlxYKlK3BZ5o2epDM9129BgmMCj0
VI6KJgKVB8/GK9dGLzhZRaT8hkT6E1QTBh94yA8O0JwQuLc1eMn+ELKK0ZZMAZyB
qNFAxWj5tQ3S06gTh9HF2wi5TP7NFlIG/uBnxOjnQC6sOQQBdryxZq86LQWPXCSM
D+kkiZRlXwQSZR/fiDxzRuf/k+Ef959vkWYEuTIxgLdc5xZshc4z4EVIUQ1BNy5u
iBsSUTid3lGgVIb1K9Sol81MyREVQiLyTPpEABIe8sZKIpevjF7dFg6zR1NYW9Ch
tOfAc9mIVxg48mapS44weDf7NDaq5OC5UvXTmxC0YqwC2hAxZzscwuWhm6wrswNj
zHU0AYiArJ+ax3FGoLZtoSBl8Y8IsPLtQCUpd7uTFDI0CqSiNTVszgohM2tfDtG6
oYkj+IBxWs5RhNuWv57ivmeNXtjDjIv0E8EW2v0jCNhY9PkPXpa8g6p8nkO9enmp
0TUz/a5JYqy3BnCD5OfnIs/dAl7+NVdS0qNDNz+NZMjeNk/jxW78o6YWMybOWFpE
zNFNs5fX/OJoGaLthKbSYOVLXy1OxMLWtod5PrPGOEdj5Qf/fQcZmDt+WIfXzP8W
JiwDtn09Y6dEWuNbDoq0l0q2B0e7BABmngC3O9TVTjiAkF9LxnGhx0f40LXovVGh
lvcQsF06h8NOeSUEsFYQ2DeG9rlRQTAMmw3eBUhMhJiMfSlZVN+7eHrTAzLbtFcC
nuzhAjcEdZErLthirC2Ubrh0VP9sPY6Ll5w2KlKilMrh00X164iXnTxnxn16W4Lz
K92YEPLT9UchAyVEUoWYnbyUj0nKLXdKlGKOsrsEJMnHxf1W4XxVqSOAXbol6JXT
rOhflwuhiuLxjQvYbrFD1f5086xkDYd2uIOYIzruhQO0Lb9LPAL6PX3E9uYVc6XQ
zXop1A6trPJYptTf61+TbXKwGyCXzMyV//kLDwM3Eu19AAPsi7+uVV2AsKlc3zaj
eOyLQKKj3fd6mU6v936R31drf65E2XnjDaEKYaJ8i7k7HdaPjrH91bbM79Xql+qy
7MyjMZ4zkIPYlK4aqrl8/9S7ibQRwsvLRCaKlX5ey8b/Y/AxFPe7tm3MpJGwqUGA
Tm0cH+kElE6n3Vo9lKuVfRNOawzdEpUYz4rJ/1/WRraXXGU3SpHPnlzO+6jMkxru
B+H/17asEqxMAZ7j/GYGAmvi9ExgJZbqOgQTFV3fB5gw6/ysH+BgDmxihpvXZSLc
LB4AtmQoNkeqUOO9eWrCJOZdh8et7tjEkbsdgadEBJ1Pj9tBiFYS9rpR+7n7cHPa
xFgSgGAvMJH0qQ7cgbvCwJZWdrqqIFpy/ZdsbxyR6Ox2sdYe0w7oFSiRSXWdqPC1
GVtsPQR55Z40+4r9/koYrural6pqI5dRnaxjeVy3M7K6UMsmWFtXP+RqT2YaBTqL
pLcrPYfJBaiPWIBleAjxcoCNxqYeAT8MNsnNvBpA8AP5tujYTznu81NIEVrSuC0V
7bhVsIU7gP+iPCUr6Y+WIL6oaMgjtSp87IZ3iMRCXEkwflWZp1AZ//NBtvJAFSFJ
Yf0FXDyP05xQ0RJ4cF/tkbtPgt4Th+KfUJScqD9jXwN59mLoV6QtnypDicgLKyYu
0bLamoZ5E7mYhowtXhlvEQjex5zk/7eDKAJCdXTUqEtQI85M8XJ8oDndM7tn347K
oGu9K0zwrruS1eyxRyc166No6vi9IvimR+V2m2pOuo3SeaFApQj9BH0finiaxe3O
At2xu0DEpDT4IGzAiLWYfvCOWzXf7bjmg+HM0VxdOP1+Xvi6gIazV7sl6HQn4ofR
wtTn+ew+gJxlRnmpKXHSfZq/g9CU8McdMD2de49B0s1/a+2+LwTahU9GOrpRj9OX
/5D3m4wNalO+5JFzcdnfIHqpDS23qmpjxyvXWQUTr8oJ5s7BGv2u0QAcRg2NHOJU
OVFNwlYwy41SPXm6jNtNw3yDvDpCbA64hDJGbW7OkynRubzclEtMuuDqXAwCFNqN
3mbF5ssFCZv1wRcUb0mj2AgJWmNncMHZURCMJlezctW98AvYWjl/hRm2Qw4PQ3IN
VgjoxrjuitS4j9/oLzUErkstnMv9F1Sta1/P3HrQH171+5gfOIsQLkZZN37gRrg9
hgRg9FC2sjYgeoGTbDyMBup9gCOC+o/m29FmyfeqmZ6hljpphrstHAInzCLctX4W
rcsDjEN0KCm43rYc9124kqsqJ71PQSNYdVXO8Gjhtl18FvNPt8kABmBHf5XzD/J5
vUulN0lRn0Xpqi60cl1LISANDD1ovtHSSGOOfjXhRe9tq/yTONSYUmxlwjvlxzv7
mPLL5mIwOWArbmgbtMdh2ZSxO/5dP9//axZ+7nECvVnAAKDktUHqaZoxjB1AP9Fg
0ig+ErtJVAb3nBTdt1r91qHxZ6+mk+lOg47SqxwJ+hG4KNhhp9L5+YP93uqhDVBN
YjBhABuSd4geN1aR152b+q3SLPTNyobEW4D5kheLFmDwlt0XWa2eEA+Jq7TN0WJ7
fHE8hG0yNY1YaG7eY5FkLEdi1wieSZD0IXqBamBSNNRguHF7u+O1FlDnUjWNzkdM
7+FigVCUjDKXFbEQKKw4YyYx0nxD+c+dfOc6PjbetQ54SWu9EMgp37R2qFjDSb6e
gj01zToEIeQcD30YXySISEiUAH4lMTR0SoJ1iHQsIn2Tr6zrZIkCq6e8MWiV8ASB
70ExkK/tp6G5MlwmoaaK6N0OaG228T9QNlMjwf+xSdQBTDQwUai5clRcfaBttpIB
Gh+rpLH+ArOex3T2Lg1mhrPOZHwu/KiOGMsj3/EvQmuUTrqhZ7g0R9oLokShMQRB
yWX92pWI9Dj28xvHj+YWfJ36xBhj1i9fcI6sTTuLrKrpoZVNgdPhBcsCnYcykKWz
D60NzS3Ex62ul1+Y2nt/4qTQ/41xO+acYihMcZ/Z5J12OOScagoV6VuOmmtk2hXf
YEJKFhKv06OR3vvr1xoJp8S3yMSEm3LDA5wheyEcytUqpQ2BRUP7FMt0+emceA5B
mF54WaKWqdccNAh3xRGhtkPaIXjU1oPpyIbPAKHdpYuxlU+a4lTmPuycNDEX/DpW
Neu3FZPsKnD+vneRNBoM/yGfIdZfq03J/c6sgfeanaSDw2iQTTzkiJuEuK1Y+ZZU
XbLInI48A+MiiHMaSFcd70tE8A+JMxIFl5A+QYUrnCsUKqWjP9HVrKWn4YOOKMkD
9Z8971x0bU1kQJ9PKraKmkzVz4QFCFDYaJfZO84PDSGPoWHoe3IVtZCQyyULydE+
VJIHZs0wstgBKOIUl7ojsBUWjyMKDEoffeQWyGa42b8bbExhvw6yX8nDVePZ0FM8
h5wH6nf2mvfpQDbdFBDvftdJJBPcG1s2sjHOZMp69iEBG/vqa1wMF3xzBzxZnQCh
xc0vcZllsXg4OJ20AR5KbLh+hR6sYrMSkC+uWcF1jvy+w8qxaXttuE5V2+RXjaEe
PZpTZ+pgvdWlc/H+2QPoAd8E2fKXuANK3Ip3EmiuSUqJkRaZkXpdTCpOBKT3fUyT
n5RFDFhccQKT1lKkT3XLl6CUj/dQml53RXhmTi2lIyUXE2dWuOdXwTxNT8a6MyC2
3jM+rHy/Gc432yYlpmyv2/BG/NRM7A/BCw+AWFaoMI8c94XrtErmDGzWxjT4ohQw
7EpyKjXbMIzCEu/ZV6G/6+c/zjnIBeF50XJq/veMYdrzE884IMu8n+4z7MAMrDYD
dhIStPuFP8VxeMok9/P1wTAgGS+c6iWtNXvcbZITweH3Blnyg5GccU17arodyIAi
v6e38PTXh8qY8dvYuhuG/wAuqe422oczz4jyIOpv72QgqGMwE4cncJnxaWOLKCNT
Pl2056QWN42sIpw4yksmly2BlCMmYB1iu3UkCeTrEMmxbaeTagn+Ht2Dp9jQoKHR
ciZufJ00zvIonLDbb8Aryq/MdLgFyTbIjmaYF0rSvlm2wl/gqXp6iRTuzVQP7UGQ
VBPnQHE/N4vlxV4tFgWy7ua3hX+Zdl6n8wA3XKSCyIOQ/4ZZnYVJ/96qvPuBRJ1p
3oXXUwPDX+umWvUYZk49vLt0umFvTxB501+8CNtRqV247+FCzhZ1PqN8Y0tCMa2v
jSxt+uoFxCK842vJZgNuWAPY3n6+uej2kMANXr44tQJOJUF1GAKW8pGrioTp8Bzk
JcoSUt2GsHaJuWGJ8SPMhzCJQcaiFrz11n9vDfaRYzcUvOX02Yn6tIPPVzdqBPQL
O7qUJ+GoDFJvDQTii19KimmfCogGjqIp1WZUYImea/s8c+t8L9VVF2j1dgK8ky3w
EdvS4NXa161A6hlDyM2HadZ04XXgt21L867GC256qYteQzi6RMvS1YJp4BGHyZnv
9TheDANu/rLvuNevPwE5NTIHD4VZQizmfKMqIaWWgRh3MG5tOfSfNEDwIBOEDMZe
uxPtpTFWIPfuIXzEb8PAXTc2vEsNfkh8lwesnl1TYPgI9ludEh/09hSema33tAhO
wKD23VKSC4mPitfP0KVKCPoosuzy1fGpTMuEQacktaHiYPKHE/6Z0A3bI8AtoiBn
YbPL/7kcQqhfZ2+nlI61oguawz/07o7ZHtzAm6XGZh4MQXXdIBMtgQ3zthXaXFsN
8VaHJDpORrDGXxqtHCi6YPd6UvxLaZ1bKhKo2/7bBF4Moo+rPIhX86homkhiIMFz
B734aBvMCB5JCMibEWkq3JiPWUB05F5rKiMIqpObKYPNa6XApkpGLKpKn2q3kFLb
XTCG7i/QYMsLELFEzW+9KfdZJUJc1MLG67RH8+pp2UIWBUlIjnPYMe6uHvdiR7ag
raAyZHDAEYubwIvaromtA4CCwotiyBe7GmJnsjQF9lqRDoFbfQH8fwxLB0YvrWx2
BNFimoIakDV/vvfjQCxs+n5BFfZdbPtbr2xyYclfB1+uRf9vo5m5pPnhvDVfm46h
NyEbLBveZpvzbn73hIKZ2JBgV64eVqxd9x2ikQSW2FM3AV+QTp5SV59kmwgwmSYU
vopby7QSnq6k5INVftrb6LIYv/dGVlVOCk7/HLQbo3jeu/fz0cN2nOCYNnrCOHyl
`pragma protect end_protected
