// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:26:03 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GVPXqpLav+sQolRXZlB/eL3jjOJsFK2uHtfgNZjOZNWRI+//ZpZjILEJLNAnhLKL
wwvDCXU5bqHaf8SCcFsQ06BCuNfvx55Ba+NiezATRl110aVkzfZO7OBDn5DcRE48
Lm2KOT1XkcbzvlxJgGA7n6hU/96b4u0iRJCGBvWODaA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12960)
urB2E0pEf1ZALQT7WNrduobtxiGWG1l9qTKNXyN87BK8qN1yy4qJLRC7h1+V6U6K
iAlhQUPId1oTBXRVILl9GrevV5+uJMWcwzmFDSJi7+XlBZIVlBhcHUK3lrDG5ETt
Mv40CRiTJeQCKMJzRauKE3v2IGf4L6Pcq5cYFKHhuZrICeObsxbEKVjbJVr9b18B
n73xkAD/WdlZT+FPF175nuSQnDG9/xSnj1AvgAO4py/yRLyRlIPHit3WdvZFA/nD
o+dE5TmGA1fVUL88JOYRoRnnJ2q5La83us+cAJ1+Ugqu+CmM8xyZCqd6MIYwBTay
aBl/5vsaw9TyEgbTrspKB37/unYak9hy2C1ihlPfHfIXRIyT5fGqwxeDVMzXOwXW
mOK4IxgJF0KCBpg3eFuMF7tXoXKf51JBM8YGePB+VT9G7W5Jzd0cWRXjyKuyiE4o
93zkW9eHaHM1WkYnUrV9PuuebTBjMFbihkpWpS1HqZ8pFp1KdBNOrJBFJjdfng/P
zVc5vMRNbKCb0Qoycx8rlQotQneG1xOxJYhbgNWLLGZgPzvz2VjFyJYvLb1b9KWU
yJXunafGG/oi6+Y4X7+xSRhERcG5PcJ1pre0NrTwb/QK9K3GQXbbt/yKGfkIB/oY
oMMZ305jROP4I4/i2anO+vn78MyStJhVbP8x/FOA04a25qOjCpuhARTXnVdKjsmg
mqXpHWjQqhjWtvjv02FQzf5T5NBjb9d04feGz+xMIjzyoTqDxCBzWYaDmJvCdGXb
yJOVnXZsFU6zSQ4Hsi+gCbZc8r76A7ahdDLnfW+/H+2Di0eIAFPyZFTrDPnXwegf
eFTiUoFEw+VLPpPdXa1jmd8FOU5AICxer6QUF4jTcYVBxvVrAiSo2vEBma6f5Xyj
DLZ372QMpChil8TjEH/qoUJeQnU/osO98nVLJXP/Aw/L5wsGcnUJ5hwF/OrBRM8y
C7cn8zvjGWwk/jamSH4HAnzoJzsR/D/hxkk7EZKrTpP7z+XCdnTk6C1MrxsJBlZp
bRSyHPOS9+D0vnU6T23cKviYuqIXAAFTHUsA6o4SiARv912P9hwa9xaO601seBkz
2FXvLyGYt4ssxCUdkFdWCh3+gci9/hLLSsIGQyFWIW/sOWLn495m9L4TmS1My1gg
ndn8VN/0NNbDWz7bBD/n87bTuJ5wqthqxo1IXRbQ+93SDrvbOMR89Pznjv2bs8ax
de8BhUr8rET2koIdE2xdAX1zAFP71Fcj4j42aNsmDjua0fkPgUOyN0m73aX8Mcuj
ksbbA8vzc11kdBC2wA61n9EGdTb+lPHKsIase46Oq6MM1pLgYwJM5Al/XfeOTLc/
GoFvAWdfPJ2+eMJlQdgiNgrYYqs7fVcVnQ7u5hqeNymIk0bfkMT+Xga83/Y08rUS
pk4HJFCQ3crxa3dZDuweTaAVbbel+L4+qx+QCy98BgNvwbpPMQwcm5VgQQmLlhpF
HUBsiM2SFwVYVqOKSMbELC/3XhY164S7WAnfpsGJplXjStoPlxczdvnX36aDZrWX
zmR6jKeyYxWV6cxeP4Jvz90s5NLgKUssdIzFQ7y27OiI8ndlPbc6YXEWbJ8pWrZ4
HuSlf0dOXrZTxtdEix7etpcLg4KicacV3ROl5XebvKObO2Ma05YiYfwWZfU+mbZC
yAZCYH8hYY+KF0FxHv68E9UgqPwvmuGRy1O87/g8lWDdQLYQMmfdW+Cu/a6KBMfp
lQHlLrGGHs88aBWFqyX4GoCDX/GSH56A62ls7BLE9pvVjK3FjRMaFUuG7tUfo52p
CHkAxtSjo3yFRT07Hp9Vstk+yh0QzNgewc7fSaovd4Jac1Q3fLuIhUqnb59Q6ja/
YiMNmhx9xNm6tOdz/Rir9+bttgn8G/E2dwbtfXC3p/i4JFbX5UawNreuS68Y+c0y
qEouSEpnuLjHRgjWuJW/STU+U4CB4do6BEA+JgW5dlH1rZ64nHWXwh7MZGnS8JM5
4G/mHZcJ8DoPtME7XCJQ40T1Hy2JNK/xZ1IU6dedE/cNrCXwyLSCNYXqhV1eupFZ
E/hf0l63x6CW/FWb1F+Kp6l3qi4YCbjNE1vm/brXhFIHIzZEFzJjr+t5j/qNEhNc
N6QMyFROAk8ndl4SWK78VINdPE5QNhsqvbVfd8NH5x/nHAXIiWBgqzrjI+4iB5tg
c5aTYqiYlNb5wEXMo8ELfP96thdkZZUyh6Bdby207CHMxyqqqTE803vn7QFwjImA
Esm+w6AIgXH+oQsNOLsbujkXfeCZH3pPGyX4tfoy0cH5lDbqKm+zX39DYnQFIZnO
OQixoL//iXZvrLVWKs+/ybVoUgH3aDs/h4onKxDjOMifX71p1GgIO8LhnagrFJXS
AbIxXlsLIwbrq7aPXUuRqv/pp+X62oUugaE9dyPFj9kCr7fJUBRGDcjhvQzVYSry
/OxHLnZLCtqiTnbw4yKWITThuBrP5idpDQX37BFOTxS+KS6bYCeHse1BERAWAcaB
mbLppY1DK5dh9wAujb6D+3iPqdaLdnM6FAxqnuZyS7pNJntZaRf6qF+Owh7sWY4K
NGi2seUmj45x5pHrzMpvV108GywEwDrEbgQMs8cuA4MNbTumek03++6boySVgV29
TnwXu2LoMs/lEbRkVqO/i45QympER4I3qaF6lKbMLVFzhJvX8kpf6JXrJt2kj2fc
27Gg0TbP9cmxHYI87sX/GbSXdIIr4B5MMhnNqJdKXd3gsu3qkuvaDL5wMGdayllr
lATRiwAVshqhNQPkxMtyc9Bj+Tsecj9JkkABOWpwQPO4B2yggtGV8TbmOj745i1h
6JJewTwCbfDa2wLTZmSoYte1VyVbOQM/GfX8WzOqAK52YUZS55ztUkfiJTKK7+jA
awOJ9gZouTPN4dh0Yq6PhrUfC+V2u0XcmK49TZGvSPbId6F7NoSW03CaNZf9bVH/
jomivQwl3icssUGxYPRy13zJQ/OzSGFC97YvBNNPi0fbpP4FhMjv/GTvbymafQwv
2B+KG3pfakieNbhgk/lEljlRibOLs3JvrgoJAqyS6tT73L2ieJq3ygo4Bp/xzF78
7iDyxKxX6ElOfZMerpZR+6DmibQchtBPGMeO/C4Jzor4L2pV9I1xi/y5s7+ZbOV9
RjefZfZ4cPeix9qyUVMh6CItpMY1Gmsw3G6UTsWaZDBYAXNCAUoj44oywfb9Spsl
pJTdpe8Vd+MOWySBdYWqL6YvPJt0HiYlpmc82W7QK3x0RvRCjSvtFzgJeO4zJI2H
j8jup7Q260pr71fEhf65H+Q9djlSJLMNLhN4q59hXwbbKnfJ/MZe7bylZgOoi4Mj
Xk7+Rob/N/g84TskJsUpnqYDCK3KqZ4XVlgnr2wk9n75IYjOmVAusn13ENf5fA4Z
3jAhEgEpSkQ1eVtDQbHyHp2jqKn45WbSlaOfyxMJBVr3eqKzXlBpedHTL6lBV0+3
WwwDGHZCWDL54SbQyua0dzq/IIdtEc+upYD8fi0v5lac2FUCLxN8zsdA1G6Cgkfh
BPuwsqH1wadw1onXfrhGFMmYdkzo2aP5ZBlog+9EY/Xq+69OrADhNu8YBgguVIUm
mKDDt2uMl0w/g3Az5si6dWvRtTs2OUANezFOGxArHWM25HgvChmlKiF1AtL4y8G1
kHKjuSfIdlBZglT7cF2fJhsZktmkVJe0kfFFUh0mscBIKrEWQFeOoHzN/255PtXW
KTrzhNm7cASp1gGfukUKTB2XwK+oNxb79e4MLUoyW/IUX/woE7fJw0UQ3iB6MPzr
fXoMJFVnww1ToOeIQ11Ygomc4gq29rBK5FbZMIlEieLWQqZjXC96mqvRY79jOf+G
NxdUvD2DpTGhmTdbqXs4ohgy+VH5c6L5tgyQtUAEnJWTuf3fLg9IEvKyuv9sN+18
kuwQPKK1XmgUE71RtxfuDttyqDAsbxDfbhqNEiNK/BgSm1aR1ky1rIWwAHPASUFy
3LYgpAvj9odpRzrhcLdLRsEj42GbxJ8SEQyfLjohdKR3kmB3J4UJi61cEf5GQXTd
oE+39yixwJQtkNipAscCy0e95JNSNggNAzSjJInaw3jWnXeqlJH6bsFlhEYQh4Mg
ShIei4KEmr15d+TTkK9E1Dd1bOngxG6aKUBVtNQXnKA+sgShFI0wSoEcmfiawm+T
Z8lgT215aU3VGRchtwlXtDMhNdFtDM0p7QmPvJT1SpiQPZ4pLIwWJoBgyY1+Aqin
vhPDYvgoCq2q+3zVZYgMvohbvFsLF6Ko7eUwzrQ1sLt5j/LLW/zQTwFRZlfNUZPH
t2CNE7W8EaYRwYFL4OEfmI2ORUn1aktz7Wq6QbEbxG4pqFJQfZon2hWtPjHw+yht
63quqpsTD2+BWmMt0JeAjDp6uBmd5FvuLLWBzumnrTNsMgy5U2AA7IkQRHmYJIYb
wsOOd5O0kzXEl2h3hAVpZ6h+jeR9fwQxfJf/9wx/jkA84atAi487PWkBe8y2cqjH
XPNf8l7AxOQm5+cRGp2LgWCusSreEQ5ljpNU+7MCOgDij1Ketd7EmwcR9Cm1pJH7
rwjmqy5gvyxPc/J1ZiwvXxPNB35FjZszc6qGoEuzgIhJ19OhdO/n3BHIIIuJGTpZ
RQz7qumWjoctgtmDq9JaTyY0IO81n/l1OaM9MrcgylfmojYOfUDtKelSyACLhwyd
fgNaNMLM3ENEn6koEMKp4NodenNmfOcKbUIZNLyvq5lt7dR807vUwI/AxASG6YrF
rlguzFPYAOoJ2RtATC5OiiA+WjqGi5MbsXBEWkFwXp4zXCV/FAgw65CjundXrix4
XQTuvRf6jPjHvxIqR0uNrpD7xGqcbQJOE8chEmgNyykcFO842esnHQxEShl8ZYdF
4NK4U45HQRff0j68Lq1CcFgotOqc2xujVyEY3pGpggggYHRAb9X8mBMzFhA25UQP
xCJOVuRKI0RqonudTnHJPJCS4uDSdQ9CSEi+AOvfkxV3fdzTh9ZeQTkAmBbLCo6K
48Cy3175I7mkYu1IWdqjaUKxRODkci+yF8x411+RKbb3iUj5VQHo6urIlJatT8d/
W/+k9DLaPntKNf5s1E/s66g95Z5MgXHcRyofy8zisuW6yhPoixrJ+2TlU9My55A9
CuY+70DuljvFeY12IzcuDXVLDjre7rIrux2/hxdwcridVRgu4fCy5T6HYsdpK+Fe
XRGnYmvyRAj989s+WNessIu+Vs7X6GHLDRnfAduOG8p0JulaslgWk/L1fQMKP9XA
hkXC1o8sI93YjhMotgsVmzB9w5w9/gCxnrCWgM9EQT9DIquPR7CBwODh4/E9iYgc
s72gzdaRjONpTY9W/7Lw6XtCwQCEhniD9MYYaS3d9jHuejDzEpp1kaVipfLAmiV2
8JsC+7RBujjBeutVkgx2MnhXx4En2/hAaGTEtAB/r9BH4HxBCdv9KXTOguqSs4+d
oHaIhEUsK4WzSAYmAOW8/Z1t+wtJG9HBp58c62TcCzm5C69sretP8/rESvwmd7uo
GQvGWeOyf0ZaTDQKDjUN8FfVoPnD4tTCCgL5KZd28399Ox7XGdTr0Ao5VeBettTh
cujwrGgCNpFd0uX6Rcg9xYxWOGz6BQg1vFKRI+7Lfyz4iCrMQ6dT/35/eJV14AtH
G6ymyouN8w8Vyf36T2LKhOW3PzMZYa7LcVPGj2bqDV2l9y3eWPjI4K9BA+YoZb4c
ggLlOO8bJeQOAY6teUcrnnKlJzeZe/mZi0TLun6QK2EnYAU9tkNPnkUfeyG0IwGP
cIRA1cLi17maL2jUc+Y2s/1wakT56MNuPVirZpiG4Pdgo5Q4IaIaWjYAXx6UAXub
VOFbDpdlQloehQEfr2AlzRB0ucTOyxi60YO7ShrBpxpetlHq70RgFYjMtYHuE1pY
VFv72VWie4bhmybZaCky9j4TGcY3kYMiENzENvjRfwAITLphlbW2NT1jgGbCh0nQ
Wq0wSr3Iu3CPeQKhOFC4Zn2tiZ8EN6BHRr8w1cncdtW16QGVyGHvQj3S11MmIdmH
g8Eox43zy/UBNBB8SturhB0fogzsSQWtzMre/U6sPH6b6OzKSjctiBJonrX+tElq
SUL11cOqWIeMysdnkb+HRLYbdUcYfxNyazyOicwEYeUVJYu3REeB/u8C3XXu+ETq
wg8ghUSNeA9+RmqSSVbDZWD6S3jbOjBgYnSCmWjPfLLttMHbf+YqihbLue36N86v
RxG95pVz9iUSXb4ZcsGmo57APMvGgtB8o59U8kqCSIpvKfqkW1332NjiEey5atGT
BprJdYFeN+ZSjhfcIOaVzGRa+g2ssOTGgXps7C+O53C4ZC5Ys5NlkWQscB7773X0
IdRMNkrM0aRPJLEWQlL2gDR96UP6yLcUIam6phhvd0N8hzKeZfkOu+LvdMc38n7Z
scck/Ik9r+jQ0O/50GpzngUz7m8LKlNSy9g6ZM+bs/NLWZ0xjeICGWiABGf6NfdF
qO206h4J/6awIJIpUjpX5dVluGxFJcCAFLTkou0A1+d6KSIbJnDSUIkPIKAfXaGu
g/B+Jb+tuyQ3nSwVZSDib5E+1CLrKdw9IL42MQ2iLiR6IGDzmzPiBvWFC6xR3Qon
VzkA+e3Jx9cFJkijtRZzYCdPnzWgFxhuuXqZ9zKiQFwDTXaqwCq2vSgcI/Kw4jh6
BoHTCSBo0zHBiOknV6fRB0fLmHcjatQ2sH00Oeza+cSTbBBbgSg+k+qNVLuuxx/A
ydGP8OQv9oA+sLfwBnF0yURhYEA5vrcxICipGjMvjVbdHzhg2t8iW+CLdWy9OwhP
qb0aQ4bWXYxQOZEV4XniB0wXmm3mAvzrwcqCDPKgNDuqLDY2LM5poE/LZVOKLeJy
T7aALgbPh5PWZGffZ4pKwYM9myQL3l+a9cpG3j0cdtuZNtyCnMLWTcjW2Wu1eoEI
Gr9E2dLIo1tgTScPCxyyyJ0h14r3xvTVU1NIguQsL3PbYaURJ/7XQ2cZ/xcLmoKh
gDcZxVFtaoY0puTxQOF2NGBusAPajcAaOqwu5byxaNcHSP9DaVCK1iTZIvsyyBhu
E4vybRiX7xrhu1PT0/oKl+cTuvBwtsTv09ghGWLyF5nG/3IdY1EkHO1QELOGfcOy
zzuLdyulVubczcf2xtRV4in3B0xz8rxprnpplHcP9/HQF0lp0NzgeKB6FXHpKgtq
bkJUTp0lndpX7v8i6uetGQ4WDLDyqcam+CZcRBY3K6HgNcKd7DxT6FKHhZlvu4bc
5WwA7X0bprfjb+QC1aa6ermOnRePhcd3BeJFKa6/gPFAF6FKM4yGK4P6xIbYLpKb
D2Ty5OVitnQzN6n6EX5h223C6IZLODBEzqK/2y2Iwk5+KD4OKgQu38rrFTaKeM1z
4b8kV0SuLFUt89STWEfKbZ18e5JXyorqld9qbMXGTIFHzqitK5fW17mt07Nvyotw
d5sSBdjW5jhdlK6cvlD/UNj9Z2ftEsbaJBAWX2qoIwaAMGNwmT6QhyfR+aAbeotH
z1eFwJbjK96XRXketv5IgcDDFRlg9TxjnyMXXgcLOS4I0H45OY0xTrc+jmWQV5Nj
gv3CJ7gZ68OOc1BOwKl4bNaUxNv8UFSS3pm2BILu6kj6GLfqDOCwf88lB2wPD2GF
vt13VixY9i28SfIznhwkjxVNaY1pA1stpdeZY2GnlMjiucfNfqZZeXMhXTabgoCb
2h9tYRmIAZw1iaNx4MHKkDMPFDtaDIiTfwaAfH7Hc1DdpCTYXbWv3pei0yBIFH2p
H+uCkH0Rk+cmlR0a3r4EsdjgmzIjVzCy6iv0sLoxIcoECCCy1jWvdf8kkrFHn58m
NNGvPRaitmXqkuvRgz3iuChFmiZr50jzIm/9yeV+bF+jvlUv1uECAVlwthxe5WQl
JYnhKg7zZWgK4VKcRUXFTsoHUqXSAJmMNqX4i9be6nGlPGyLFcQfniY5B1m1Y6p7
EtZdNryNr3504uRywyTNP3auEPzsKSpIKDTl0OKrAtlDBsKmU3/zO3qZDcaC7ZBT
rjDUebzXfBkfp+YSxCAUB3SlBWSR+ErguZbVFH2rzwA9AqXmyrFXAq0sLPy262tB
Q157PdHatlfVQ/DaEEnRopfRW7iATexUYxDWQSJF1xAGKAmw15tsosKbH+AOPitz
BXaNgEKHnGABn31unhd3kI+aFk+ZirKyPj9MWyVW+xCWst8uVw2kvqYFWXbAbdDm
B7XBbxcLCEVt9xbY83aAuGu9KscbrMtm7XbyNtAjstRn9W92NjddZIHD2mT3imXG
tvxflHshlOqLzLcBHQqe25CrsG5ELU7ldsvm+nv84pdetCJ9anRUGBR2wfBlWiJe
RdhYTZtqVs65/G0JrlEWEFxiteknxzXImFw8NODzNbNjHiAp/ISyjTQfFZrJG8FC
Im3febmz/v2SZqPKWihJpBGyoW4tgzbY8ZAb5Xrqrhvy+tcjAiDrSS4QKjo+zdKR
YQ2BLrANlLeWUmH3lskiGpRTqBLT8IesD9QSTcZB3eIBVRAV6V13TD3dTHfGIddM
R6QvE8LatID7DleJZRG8Eo/gB+CNYlG0X7zMZRPXlHzl+P2ZFdJ6dej3VI2irS8g
cOM8ukhATFbE99Pk7h8vXyn3EDsDbGvQA8ZW3C4D2WvqxmDpCSs+zs5T2JCzFDpl
L+/Tl/eOcQR3rpfeGRU/OC0+uN0HoeAaL5sYC/OlCRaNOET2I4QxT3gTSTraLSRF
vXXZqbJodi7ZnBiljohNfYCSkV/meInTSmNCjZbSVBwlK6YHwxkLU29DyleW1a2O
SF9vkJLVPI6qv7xN7QeJtp1Fm2QPxAkiIlXgauuYbHJmHSWeWpfMnvXGMU9p0VR2
0RHPGpHMQSwRYJunmqHRt+PWKxj1KBoBOBNyokCyLFxwLm9j+afFba4e4FEOoH5p
JeOnxAipQcrrDZ63psSC8/3qzF5Ndu5C37yY0b6eOL2T2KtQ8GaxueCC+Jje/Um3
+HJ+IlawDRV5/Klwy6JRQ7BG137hUtOxP4PKzmMDkeYLMcA0EdiYkWdN4B7stb7F
ShqO+eMY8WZjZNP4pKJ1yXWgF/BBGp3ZeTgYEv1GlS9Nc9ZPLMdsDtzkhnlCZyMm
YLnPCdwGUlsFFt2Vi+SVzRgWqtXCJ890me/fIVJexc7jVb+sLC6ishDknuQ+A1zS
7NZZwXj8EiSjRym4jEtVLVbPKHSLt9o5ZT/6EtQD5K/UhH1Uy1fSumXKJuXyfTz0
82vYxIj3gb1aEKB924REzqScD9RXCwIel3KiHqL7cdG6z2xA+GYfaWCTMDEXnSEA
BtVKaj52uXngGBfmkIVIyyh+QMft+zEZOgeMDY8uM0YWQEoWt452ggINWlXY6E9P
i6GQQfDZSiPSPW3wSpflKRvCqEaH1PJwzFhqJaFzUOcdYL24W8J8+bx4sscnQnwD
yQV06ax37N09FFz/PSvAEnCdNQFd+iJIoq8lPlLnCFNIpZuUvfACxUqC9h+KidD7
XGw6N5MB0NG5yo+8p5Lt3GEro0nNndDzvgro7TbLS687ONeR2cmT0wz4n2/kZ2vJ
nq1yWzKcPSzxwb1oTEv++CKc+Nc3TIVWmAzNSqpm+enudiYWmcU4aTFfqWJ30n9Y
aT1hlif+5rYZsnamkivRfl3AUBy964ucTAraC9qp7OEnjePPbY6guJ5n1VAMnk72
F1GVk63v2WQGv3dAv7IKKikDse0IlONGB+rHrjnxake7P52ojgwHCMMM+j8x1E33
Z1dE1wBIEpl/Hxn7wCfwkub44pPYeVxB/eY3B5Tvw057m1idPKgmruCcFoCewcJ5
igN+QhZ9QT+YWa/ynVtVyjAdAq6pdg8KKSuJEggDppBgmKeDNAlhST72JUVcBZOt
z/mpWswNjyvLjmztg2qN/XFq+AEvXSndhMb4z4lKsm53XP0dJe+lLAaHbQVm+/aa
+KgMtj7XjCiXBSzJ9qUqLUBkYQFfTE0c81+RwUvu58DajfkgpH+xC1yids9yIj/f
Gdvl3uiOfqQPwX7I6msgVsSDAjj9F6EbVC961fbKQpPObI7Czn74ky2XMi1cACae
5P2DJyNHe4EQID9KvPI/OgLg+eyYD8wmZx0Zev9lPKGUa/NFyqUmeejqxdGkV/Zy
Sfz6+VKN0Ospx7+iUCuO7jAjYZ6q9Dv/eXtbIJN25vx333AgcAbAFa4YG49POZ6n
84aEy3XqCyQWtVpQynoh5S9ze5DxzUsLeuZXgTIktvjG7+VL/YTqDct9MKTWFVxV
2v6o8Xo6eWQ3xsgH2lzQAu/96GrDBDlu5GCNge7+MvcqcGgjvKj2VNiUEfFH8DqP
0ZcApANrXoikgg/MY209V2RtH1AzuEc8/QBU/uiZ9FlK/qM78D4hiIH+5omwzDHb
/6NbFQTZ8sn7ycmO7QOzW93wrrl03kgvXhpfDEQCD45KtK12iYQU4jfqfA2QwR/P
LQR99KMb5oBlxAy1aDZDXEJb0R5cklx2sfsmkmA06CmyzVYRkLMSS0QCVsqI8L8C
S0IjvhoTqvTKjQ1iThArZN6MUaWyGkMQ32fUP3xzIM+giKsaUga+ru7vpOVsczc9
ZTi+zszlhw7DRaH94rDPwd4om9GcQLUamDTVCQxzeEHyUFDZiHICMKI28l7fEtZc
WJnYD6laufPskWMXJrvW5cDTZtxqFvO39/xkWOJY2AvGMkVj7XePyBolEfDMTlLa
BBHOpiYzkNo1LsuV6sw3aLmr/XfmU5WKzRT+V5W/letnt7xJeXTYGiT8uYk1pCQI
SbWXqvSAhDu17wtvPaDacdE8a6S5KBqNldKnDDnp4ye2fa6kuU6V3KHAg7Q1GGfQ
FuERMiZ24OW2IkA2To0Apz/heXGiOgHeyYo+EmBCr0CQs/OIsf2QRLP3sFd7ENmS
BppLWSnz4soeRHNjQxfWQjEctBh8TU66FFFmuXMUXRQqFBraNsIMym8skjti4BLZ
WU72Qxd6YsueQxzB7X9nj0TJmk/B2VutIqR/Mcu2rbEOJODc9D7Yq8SaaTgnIlCG
TQiwMM/MQ7OX/3rBKogPaKyTXbttXq4S4Er3nBYV1VA0U4GuyaXvRMCwLxb8rlIa
M6+dWR/iyHH9SrsPgIxkzdD58rVXdMOHnoI+o9T6mmt8Yp5J03HMOQU1HBpOGhVR
ZBh8n2kzC1cf55qjfApR9oqapTdEmjsCHTv+QhEvOvyLIn13qLH1wh2Z/kJf4fjj
bNT4qWxrMndPlJkgnTVCy98vb37EVrskoE572ZDQ6PlN/pgLQWCSm79S71RMP7hq
68lw9eLMJdzorQyAy9RuggKU1cwqzTdXHpRn56674yrkX6UgDsd4foa3Vb/S8pUY
2fU4CBeYV01+TCbXNA/howZ+M0NxxHcu9dqF919UuLG9bbNQqr8jnnP1aMNrFvUE
DYtH9ZmCvqiSrdvPVe2l9whEQ5CLJhFzEP0MG7elaulkZQBKE897IXmIOGpyXiI3
5eTsoOo8ydM3LGEpTqzAIjN2j+vBrFIHkv2EG3XS5RV4Y1VfXByQQX9q2QSixYju
l0ONhe7ldskqSxINDX9WDOdPd7GTZ3yxbC5rmY/NG8Sj1fCp5yDxjZsK0uTCnPlI
Uf6Gl3gd9NB8JRVQIzbWfJimfIFCw0J9p1X+Y6yI/taxWKMDNKRnYe+8r1dvlPh6
qZACi8MjyPoRxGP75mp1o67BJ/AYkBu3NX4RH26wMvEV56Gwpvpe4uhicyXerbhT
kVsOPtsQOzlDCe7zV9wSvfcG3woLDiT+JJLhoD2U7UmyKC8PX2CRR3x1uaFkAAk1
trhVoKIQMJ3KT4cT6/5XTEgvOcX5mE7UYzjiwGNRGz9AbqAFPWy869waA22xs/0K
zSFQBWFsmJ/41ajukYBk/TpO8NcX0/Jb7p/ZOKvRvY5YHIYqrkSBqtggnNB70BKT
LnD0nD/EuWLEPmWxrAPVR7ZZfR62jbP4vbDok+uuE0N44xGm1rwyvVDNdKBTXb4A
mkqCIzu/DM4MU6Dr7wWvM7i9v8hqzB35kkS/kgYAzkJKQVTF6eEv4LjN/l+pdmbS
nB24CA+NF7A/2zfGaLHv/MnTuh8yZgsbqf3+4kh2w4gFTBIcKE5eP8SGlS4+ppbA
MjiWy2uJ8zSn9YLARI3yWwDWIcHO3EA/RMlbNREfgWR+IQMptPoS358pd0T30u7Z
jR4NC02lenwNcmf2PDDbsmN3++Jw5hU+yFIHhMyMimAF842wB+sjhX+jKwCs3+ro
2CmoreZhLQkoogjJZQUz7e0jKvvpdFD8n/yslGptJro1vKTr6KGsfXorrXmcuvne
r9OtQXb/CAvdH9gGwsB7dUtreHB593fDLGVCZQ5pDK1kv7ZICDQQ3k8epCX1OcM3
Eq2LJdsvjdWJzIl5/yXGST3t8nG86E0PPzSiDcv84sBXxnx0mxPEtaD0zfQcs6Kh
heAco5M/rwF+o084kIQFy7Xf4zypcrgmokz3yiB9Goy4DFF2uLlB3aDPlm72l7Su
GZ7gABG4EfQSNE4b4tlFe/1KimiUwAjn6zEeZ6do5vHMvAmzaSA2jHYyEPzNJyTW
tsF9LFA5FdFXxjixGj3tVzmPbIsebPNLzdzLZMXjuHAzpu6Z+X7MP/a8vHzTWjAu
0c7wpGgoDe/XWfERIFIQzqadk3C45B4MWkKf6d98SfldDFa1T22XYUGXTNWm6jwb
99KpljHXNLK6gccLUxx5Ws5obw54cXUTzazsWume3DvfbuwMjemhkqXArmDcyT5u
dXrKuECMRx2tYzD6LGKftZTixTAY6tPiyZzC2w0SlsgOwlNoT4euJTSY0mIoLxoj
ejUp1GzuHnx5rvPF88fEdB/TAMn+4T6ZaqOOK1UMnBWndpYQl8RZ48MttQ6NdLOK
jx+6GiV677W/rK+fW6baHLW4+dJsnW1v95CnTj8XsTnl0jZSKD3w+n+pcy5diRm7
NePu1cXSaRwX7vdQKHvrD1qbQA19KDWDRpaeMPxRxQ/CSLEPPBzDUqJUZT6pOnO0
UPayvhs/IurhJKhBQZhLjBHdAZXNh7Vcq/nkWAsBMV6/ijSOzFYu4h5OnKtDxQIZ
GYcbvVZA6Yy5xG04hwQR1DauJmYPTdW0l9QShQY3ZJhR+CK9UzJV/HvytYgDehv3
w3NSCtYfqhUBdoAw9FN6iHn0d+aUoH1Z5A2J4TZ9HNvuAqPvbsmCq9C9ufv4+hvb
9jSqXoWogCCIKvmlQJZRlvHL4QjsA/+mn/egHPjddltNTpoK8cIi6+K49IdmKGUx
Wpyzs/D58s+lW1kaIIEe+pvOOuLThfZxS/dybXIwMUpCnmgmkgQdFs7IQ1+seRDx
ia9yWHgIqfce2ggrOWUDU+OAbuw0fQYWfRHl102P946djWmZ1ocI0sybLfm6RROs
5a/UMwOAs454glSB2yEwYVJkeVsqDW/HoEwI5bz+OPlQ4MjUgQ2KZTPDGleoxxpi
ITUIn9jRCfl3/pqu0pDRzN4fn7FepyDGvTcTNEZ+5wrJnESYFQRVGp5cVNPfmE0o
gzLEmZnPP4T6Y555j4JHq+aqdXToz9UIbkAMXBBSTcwJcfbimb8Six7V4jZj03Pa
PKe8NpBg+PdOK9DMk94yvXt/WnX8xXG5X4BBSj+hqd9dAm8RyhQH8yxJARH7sWvj
Mjb7mUL8SA7Ub3lolJHdOY6dnlPgpsHJ6A5SosqU+PQE6DccRXKZ3yj1KSyDusLa
iR3sLV188xWx2mrVvEmzgKER+FNqHbZoa1451hNFYIY3viAlLwy6L6e99XI/cp1S
YoZe9+XUjjR0AyI8xUc6BSqGqzkBeH7OzyhGTtOcrktgGSL8NI37Dl04/7r+1yfW
epn0ziqvH1ZWHNPDPbnFFVtAoiG1s0xKdDDw3/TIRGSKkSM12TsgMdmgJd92xPgI
Pr8roO80UOD9PvCNBO2JdkG4HANzRzOt8lzeewrVFcQTFuVAv9A/11E5DeSdzWuM
wUiZB6DWLtVV+Oo1JcdGjhdWq0w8Bm7kB99cMZ+fZd17CHKoyVq5W/JS7wWGe2uk
yWEEboPoLsGARwmifUFKHIIjJchcxOGSi9GNqNH34HAr5hDUUkb5zA2K7Et3OKf/
cj7AunIIFp28OlrXhNL47xsYAQvLFl1EiXK5WX05E3IkBAGDCxu8ZDV4ERAhSBi2
iDDPUCowFzHnAwP+H2IwUZiYwqwzej68nOqajnXFTF9tUeNYtgAN59ADf987xtdU
61Vdm+4O2aeoQ2FJUXAss+glnfIED78xXvMzdr7E+5kOEeoardfqsSxblGzJeMjA
61IDxNsr76xAe0hAfuV2cGbUZWBaSWDAUujDFjR9aVQ1KaiBvdDI+DB8K5UFf5+f
575yybIpb1V5+QbpCoYwf66cTFdiFc+OCjlLguGLLHQfpUzgXWv/S6UASZCEHuWQ
kAH1jmRHfsTodOVQ7izorUtaKy1HrKVF6ZPHCXURfu2paK488khIlwTRjB+f13Bb
m8AtRJmWOfFkPP1E3OfIKHMIXzJdqY6Qm5m3PrYoQJ3wJYGlhXejOfxzEBKGqJxo
IMApEjsZaQFTynNc6KLKlYAmv9ls9o1G6uhen7VulPFsHOegHkFgJ+KjZnfMGlsY
dgk5oV/6sm8zTxL6m8Y2aANtcwSvMc9N5mqs6mVASNZmOlTjfG2QgIN5o2MxUIsh
ZVhgv6Ju0kEa+XGKfN8Pt0yMO54I5AhL4WtWNL/ttaqbOvP5lq7IYiIf96BWj/BA
IWcXsODGGJ3FCTDRVgd0hzc+W1N9+FxTk4jBjeX8QJhjGZsbrj0vpTpJKfs0kMyl
GdYIS4HfBpZYnABDQ7SArh8kPGbudyU98/watkTWhhvgVrmvBQH1z2PViU9VLhuq
+PnoajtQNTD8no8GrnI5seBj5FIz2p8W4hxma5gYq3dLgqk9BTDtLTuSRfobU5p+
yQgFwKAA64huB65k1Jqmo94wtPvd+MRZ0pr9pRnKihbQik8ISHGJUFFPhpQiZ1e1
fwqTPOKSZ1O9ceSZZOlWw29JPiHLZipjUDV7SwKp0KQ9RVWMFAIszNPWExmUAbKw
FtmCX+61s4npvJUYf7TQZX3bzWsBePBWEplNfaOvdDlgv7doKad5ldP+49flb0sy
6oR6PjlxCsnDuOyDA1KkwGf+JBUFBTi+FSNaK++b0xKlYJ4EeBi3b2WzyfSnjeqK
i6jBh7P+gmcARuHcvUsqvPl7wvzSGP5BrbBa07/Z0nWRssI0dBI+4dyWLqeIF5k9
NcN7yWwabqPX3IE1wMWKafm44FCyr8co22uqM6k6jSnX8jBkHoHY2GpDSMgLxrnr
pFVil7DeVTsk7bJIwW6SiGCr371sgDv1TzPK2KWDhKCfXWFLqtXHh6LUfz8U3fRb
T8Dllovyix80c8H9PRJqUwLytmhxJkOMgzE3bJfz/bEG2+JHlt2dyoj1s1h0sF45
9GJMeEjjY6myhIDrWKWpeuf58em0/cdGK1D2zaAKD+K5Beb+25BEHqY7xgC41eoi
fhL6vmnzC+IRonTlSLkDUPOw4yYpAqixjBANs2ShNUqTkCU9PNwwELNvE5xN5Dnb
0oT/wwKUrGD2UmD6nVBMgVAdi1d08f9Gfovx+Fms7GImB3lVcSviZi9vk8xBay9H
pyXFRI6bSHn/qTfQVNboYN4KykTITG6WGHifWYn2MOWaQdJXk81///elja3KgW5M
eWScS3rlQRMYi+lAKTNIOUMiu4TlP2FS9jgDPXqPw1kYTzGLE5KaohVPHZwVYHNv
gdbBw0pWmWTl7zFABelnoOtzkDX/YhlufZc/H2OaAkQbtQzPoFKsv8SpRDnJn5uz
yAPRP9+NAaft3IhJ82sbIWz/un6KOomw+zgbEwuOgTpkDbZ1mJ+tWW1hqNc37lNF
7us0PcXqFWBt8gSu24P0EdpR0jPmS2M5U6np9mUs6BC46TgAC5xVaWN9KFpuWCFD
ZCyg7lgzeR2rhCG1PCvkHugyd6KwO9iy7z4f0DX5d2ccGlcyXbO9EbTaJfdHbNEb
WOqvJdyBERX79VSg2tOGeGPu+TZmkobNZqqFruEmM/qk6Fzs94UlnWc+lKtEv7MU
xFQRhcvqnu17J/+CPsX+oP/VrlIWrGcLJitufw3kDV3QrVnZYivr4jcihWDOBZ38
fSnFtpraoRgyMJTNUfJV2euBzBf3FFqVjFG3LDHzvLEj6eriJZ6+Gz1TZ6IoCE3X
mkWpS7RASh2tvJ4ULpATPR2PzahuHHmRHwDuhyhFsUnUUJks42O80YHKlHQwcn76
O15fFhmnJdNqADg6pE+i8MfNIYDYE4nYz6Cy3Tg+t0YNk6fEmJKG4rbg5rt3LIug
CNtuFwKpWlSmFgV3wCSx4WDZ7vrb0cLnZyPB+B8Sb2HsjHfSM54TG+GoTQAXO+Sd
Er0tgmf9aF3lYEDeozmkCStguDh4QVWVX8OQLPq8smrrpYyJwVoRw7c4dt1tX1vi
nOHcIraxsIDuzvgZLbMGBZm5sA/rFJhY6NEtVGJCavQi9Rw4pc+s3veFP3dJzcYz
rJpT/8Bt3OMxaZM3AXUWVuyuQU9IMletcV8+Zyd/HNFMVdNLJVEl15SWgfS4vcj/
vOM83m2hKyeTBHyUzOwRaiomGwedKRz5LSGJ7hO3XKKVXoWbKKd4Z5TIdSnsMOVu
9Jk68yBYnLUAw7Kv49NXJdYaWaWI0DWQ+w0n3DoW0hNkOP/C6e2ICAC74pYPsUtq
WjngYvD5GgtIuoGAvNC5xxoMupuhpGi1Ak0eBk2xO75itpNk7uWciG/Ieax7kj3P
SmjPujFfAfe7hcLGw2JRAwOjRBLabd6Z2ytiEsqTECgregkfHZdw9oIuByR7Epa6
4QQZNMdN10x4Cgq5JyQz4vbZJre1YnVhKqqrah7O+aKwvf9ccw4KkqkY7J4mcxZE
1zGSWtTR9/U7LYnhBivJtQpD5sPmLHKihqpEerR9YNUyNVpkGKRBNCXCdYS+M5Bp
Ybp+sC9EuexyIauxtOBi03v56cN47JlWCbu9kBGmGzu+gvKx6qhQ390d1Zqet2l+
7Rgz+WE/3lpdGuv6vARRCYQS4RiQHxh38P3unqHzdzwtdjS8DmrZUWXGdDbu4Vz2
Rf2JU3wzTUEHLj4u1pdKVQCRVcUtf8A6XpHZtra/+v8gYlKq+DfS9Hs4V0ejUXaK
Pn5cquQcEbOXBdVenIB/VacfkAslywWcNkyc9wEVYePM/20TVkczlcicKmlcxN9v
u0ZKBj2PYV3Ss1kZGCTYyP5mT6z0zNjy5IdXxBlOFks/QOdJRyZuWI81rRDmvpvb
`pragma protect end_protected
