// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
YvKyISv8LjZhV6DyIw3XHLyvABNDiydJxqoaNmYFjA742wZSNmXS7TQEKm7rDP+G80ckFLy8U/4s
LBazKjCBPmVJKEzLDCcuOmP1icHgOY8xjLHZu4T8EAtU5oYc+1ps3LYIAcS+QM95nO3ajL9cKr2C
i+NWKVw3XgiKsl5B+jJfs3+wZ1W8o313Q8Z0lL1y40MxhklqPkz4Ay+jiMsEhUyBXSkDZaxjjJcL
/BAB9rGOFvLkZEeNceyHDxNE5McIVXcrVOBxzLuKxLQEB+RkJo+W4LixqDmcNZlLRNo3gXvt1H1p
0WvL11E+UngsC9MSNiVS7Rvz12AKk6a4NDGR+w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 27136)
hvOedyzx5FTSKYH2KS/KesxBgUK3DPNRIsZstq0ijOozanTtAspiU/SSXoeIr3RaMNsvv1raMDOI
C5GYSzylr8fJqLsCqThNtpBw4mNm5NgqASM3nyLUfaYmMqnZvImaDb1lmYcDUOo1Wrwu7/x5yibc
Xefu94ScWvW0Ya62k1Nw8T+DkdKLRm6SiZrfZAuw1t3hx9rsHvVrDoBgUYuiHwhbUcYZBrIN3H15
CnEBR52L00pep30K/rL15nAtAe2edaDoBqWYA+lAfGzX81GLRhK5sLsVXYlJhwgq1tEnFc0avUFL
XC/x8usaNeLnZEI1apeoVWKcnmEV+9Erj3tjUribVXTR0oFNJR/khJUlqIzYTYJXaX6c1AQHRRWn
Cj+UbXC5GIcc29VxrOF0JOTALyc4KbDI91SkfEjbxiumEOE8nh/Osp2+c5jCHtCCVCHPn5VQhdY2
xASwGYFV75C98fhHELlJ3v/jC+QjqHy7bBSg9/WlV9dZIy8vyI4LxTQgb5vx1wduM7x6nQDI8X3o
sDwvb3rlX97oWwY1C7ovtV7lbbfw9LCVnRpW8XwQqOV135XdlGFayX5g2a9NZsVnh20n/uDot6ng
Aie3M663Iq0XSAfTuxwi55TRyYIhN+eil14xo4K0ZGiu14h2zRHDwIMQrkG/yF+2UdjolYKSx0II
peldQX+Ro0iRKVLwa6b4xvsdHdZqO37MJwOwklcxO7WjuwAi7Pv+JaO/xRNyMSnn1bz2xGcdX1xV
tNa8GIS80UvKYA8N9DOKvbTrd+KHSCgRpRjQcx4aXdrMpq03X40s8n4WZoc2R6+vS81IXmW171dv
4xecU2M5UqVTgNZitEdPA7z/fzKkF3Nh14WARV2yGBydn6v1qxR4w3ciexkpj2VydhRlALDYejho
aKntmhFFtyh9Y+zoij88F6jgfM+VLGM/dneQ6MTzHMP9XblCbbXSVpUQbHNTMuFgcHSuFfC5oPSO
2BD9lqbXuXJvfW8qdHp0ofqTnhidodVhU5kGci2cw0DWMWPjYNWmZ3Kdy0yvW3jo9LVTuUC4Q+zP
dCP9EoKCDqA9h+IMS0d4dLk7Ml31BDB+xjjDnFKYFLjR1LwxIS97JBuWfXt4HIGyzxhPqw0kPhPI
5nqlwrLSJVnAr7NwABWloeDdnWHRjz3yl0jwzSZg4MsN5HXx077ItOzhmeH7VfML3d/KeL0zymmP
RtISkbXCy3SRCpu4UvnoaV+qPTjsV00THvopXy+v6GGDgETB8rFMBZaOEOcM+iAE9auVHb9bHeIy
tgWQH9QmLTw590vk43bsm1niJdO147Zf7sMZq8gw0iqeyqCCGeh9vAt8kH/s2Kj47i9s0ujDafdO
PafPhXdK6WREOejjb6cPOhHYWQlBPt6Xr6cU5E56UciLulGpny96dLlJEhR7COaji85k6YPsqgXd
DObs5JvmWZEV2Bp1jobtzjEJVmpJiVE/aui/EcnZjjkAOxTjMMpBQcDEBfWFAke7Pw66bEi69iwd
DOfwmlzfroon5o84Idg33s9N23RAyJhzMin8dHbK0caGcHKM2o1L8StxREuciYnmyl/TwDA8p9Wc
rUxGbiW4tKM+exgTIO52je87fB5MXO+Df4jQu1gNXRwYD16/jF7Ew14xxtPdspfOtWPqapccHUFM
Q4gBkdd1Vj6p6w77fzBF1QgVeiF4cjPj0rPYXfBVchLY4cyR/RtVBX7cIe0XR5eistRE7RT7kPgu
U+7OeaOd7iiGzkkZ4B7MHxG1kL+po9EVZws4xdoWU1xYOEejo8aQskTphWq4RciCUcEbhNCXP6he
8W/L02ZdSggfq1A1wJp5hRojzj+JyRPmZ9UiSRChiD1VVVRTSH5FviR7TneG4LpIYCH86gaG0BRz
6fdMYX2CedUfGg+WeRWEjzlKiD0C66b5l0dEYPYLm5JW9CrZeNAMiH7n3vXMtWzaejrj1UqpR/qu
TkNCsVrczy3MCSZnCjIN9JyyXsi9M/g+F0H3NMWBbTPLL7LDzrf1jatSfBv8LZILeqaSk6v4eYxq
5co2b9zbfmpfaPthc/fkz+T7YxEYVzzlUNrpuersl6IiyoQwoh51c4Yy9c9kJLbpKb76EceEEseZ
vyA5+tOoX/L40/GZXwtITar9vWnJBSeODjIPbCqMsXCEzMHiewrFWH2YuxuY//gdDob8shLC0Smk
xYQe24F0Bt52/ZOz69nA09Tn5tUzA/lluryxxS6FeUeVTqCLr6Iag55Ml8SOCZEuWd3kVgzaIyKv
Za5YB5DAPPeXT73ihJMb+N1dm/tKOhu7wV9dkWBCYrhYI8xYnM5ZaNnze/bt9gdAFS1Tzv2vsyEP
a1ahIvQevFsbAPn625tvl17xoknELig9EE3sfR9hSqklqeE3qL9NFxqQWG0s4Bz75Xujrn8prs58
OgC+5eomO5xZQfN4XMBHLflACvmeCzYVwnG1SHuaekd8OH9s7+JAoe9EOSC8Gzobo7wXbMmoekqN
ftK+g5AufjpQ1ABRZ1N/ZWdTpUm3jfdVens6dmKUoCNIcBL6QSWZgGFAUUeen02MH2YieboVPxmJ
75KsjEosTr7YjJEMZnZktPE/GodZndH3+Rmwm3S8ufHJkqXVRRCUpW0XX/d9jfua+gaK5Yfw5hO7
zldQqJ23hvY9OhBNRKXKqTFzvvzBbwqJvI0WmB87VeOTnP1Crf1MVnGL+BYvlPacl2Fut1TqWhNh
uGgS6Z2toab4kuZzvghY9QOG/TKordWoTyb3kZf8etNNBogn0TKwXu0NZKBMAg6aLhHrWy7iqcfh
GE9cKApw/mVJjgDyQPxbdt9Yh/8UJgyw04sTRfhWqODjXposaqTFVRfGE4Y0+QfXGEXSRnXMmt/F
/9KAONo/CxhWz/HfcBW619Vi6o25+jQIvnGiJcUmwhs9FQqo+WkXB9QAnw8znjVpTuPkT7jvFY3D
rnepa2LD/x3RPITBpAH0aRVeesgTcnMVfQBYtqZccdgjrsSXeWIsr/VkwJyNpAnimb2280d1Ubhf
PyKJlnDaelZVL9fSB12vtnvR/bBJ/ikYbs7ppLBYDzsDJCRCJonkGKrJxgd+JZhJA6YyCj7Oq24w
T/KaQMMck+/iM6j8fntQsKwn0Ul9uM3U9QTZygtruuTk9KCYjRsCNf17zs/+I5XhMABsZnrvTBfm
ZrAUxwEjUhK/ZHcHeQvEDmGB4efq/L6MxfGnbk/RQs+juVN7ai7U7hejaRWARCm7dzJlx/+Y7k2o
KmlOEUE5XASEgiErW7EK4AN7bkfu4r4qVsPWlAmuv580kbD3igeQKtClX3m1LV0Lf9aSVX7h3LDu
53meTCYsyaNIyvyKDIC/uiiOCtKKjMkBu+bqRa5Zjnb7ppM3pW5XsDcu2SfM7kYLrSyibehs6Eor
nmVUC19uH0Dkxxijm8dJcOej68FXW5lFsiHBOL8XjA1+G3rusrB5O22RymVwr81YcxAmWnLkQroo
CaEimLEWiAGqPuh7iEWD2UUCzb8MZegGouqmFFsDwL1ta99qIbZLJq74+vl/WMn6auKSWQwa1ebL
D74/gEDj23d1wR122zrcnLTn4rKYXSv4YKhMo/GjbDh6XB8yugbVD1n4CyXVP6Wiic3RNeyiRCDR
2bLbywsmyOQO0ld3a8VRroOVJLz3veca4yD3zIhjRcXG0Q+DV3f0Xshb1f1MrW3T0wjhkjoJ0HFZ
kAhmVaJw4i90bGzg/o5UbjWiARf4WshLBKO0kEmBLDWrxfkJNdu/02ViuUVeMYxZQ+LRTotznVGn
7UERGpGiVOUWn+RfXlD8AI2LBYUiJMcQplsBWaIFxigv+byGQmzg4PHYYDUUY9cvxGfZF31J/h6a
wZ0f7BAoiJ18cLMOorcv+NxiCTwQzPfbZBPz0IOJLYByctmz37W4jojnkM79KtSFOXsAYbC7bWOd
p41YxJ/HDMCO2IK7sAqraCq50t7ycgOY49EZwio6t8Oo/K9inxa2ig7UmZFRNVLFTdlMjBObC4lO
DfHXe9JZCbw+HpmScM2LrJbj+LAZVh78RCcwa6CPZ/tfyBVXbXcWUREVXEgeP4lReaW+Jh0QubE/
l7lDlmvDWhZqczMgi4iy3/5icjSB3gbxhnBAv9l0yW6Do8/q0u76Z6t4OfU8+xXztKh5KKuqfP5t
iUnNvIzQXYGU0yRUKFRHj0hq834XpkzxC63jVUeI9sX5/3PInKnecH0wzuCBZtc+868T0Dvc1I5U
JyAteKwW8WCZ0o1qGGOn9WuYi5oPdq6g8OzX+gl0iUz5vs8RgoLwt24DD7WI7sEFbF/i+VivCds8
YY6zY1r0cKSJZiPwHuBDCygiQAC3wGJVwQC6Gz8LT2pE0ESLJv1YtOBqlp0hQJ0byYRiEv5/Adnn
ay2RYYsXuGTyavARjwPMM0Megb37rBSSzNlgKGPvKBVi+DCMUM+T15PfI8VORed6YsbZLZpeZ83C
VDwQXade7haT08LGhb4WkVOE8FGyerhAbXx8nELRe6C5Wtmj2VaT5TkVb0UYvspTbGyHP5xeard9
R/3UngmR5w79uuK0AxoPfAJVZEC9R0y9+510EajvobBDsWHH0G/GP/QLvpxM8Yu6Aor9lXS8bkMF
Beuw7xRmqhDlYF0lV00iLQLq3nrLcH13GNNecsty8AwfatuYIdeO/lcLr/AN1902LhA+7B2rDzPR
5b3GL/ADOPHo9Bi/LTYSbZrXfapukTqPUAGf4IpOkNMJj5tcpBJb3xGnNIMtEeHUns0f5kzFNqbd
q003AGmH928P8Pkw15S4DU7M89VG3s4/ImaSdW2kWPjfsda3E2TBdZF5MvIfowdYpsDcYwgeu1yu
Y35Ik6x5esBnZPDu5LOdUwgVF1QsCNoTmij0sZwOoStFxUhfVVgqR85JOkspThI+Hc/Ccn3aGnJR
QR81GHw7Ai8f+VQ+iuTWcaNufy7rMQ+Ghh6h6ByudPvrBeRNOMyT9ZOX65k9rGa1bkwqc9zzYONP
wgEN1d//SBdbkXPkUREhGu10mGbM/HRlVasrwYnSuUI54oaQhQXYtXbpA7MMjChk3aqMJ8XQIXOp
G9nlHaB+2VLSFxvYSGptiW2qIrJ92OsGgkdqZEW10kbHU/dI6Kn4Wak9O8+r8IrOkSiS+h7sQxG9
0NwJvXio1tWtenwhBs6saTy551FWn4IqKSK+/PqTMfX9sZAL8EKvrom9Bn5Y5M3pKcm1mMpmAhZ8
PtApZj1ceEF1L6qlb0b8q4E7FNKfwLy9QblVqdIWXCaxroCaJpaqzAFtCFmyrKnwWnO1RW8VqTIq
6Z1lIYHho6/LqlHEFzQg4+D53E22HZGYyR7dwP9jiot/7MP88lD9b+haf4P4x3ELgpYeBn8ZtSS4
iibT1UHbzFACptFvqdjxr4YyNoiXTx+dYrJrezPshPDblfRfWouidnDLQo39Pp0VL62VbDOpIj3p
xmVT+SN6v0HWxKjp6NmMo/5ENvo7HOWUfkTWrLdaPiGVKWBGAyY0sYj+CPxfpazdl7NtIs9DAtc7
7AyQVmwQE0saMYEC1YcdUTi9zYT4wBRm5BUvln0ELrzvxhESAzgJEua3zHswlxFmQ5tzCbyI8FGC
IBJCcP4eC8Knhntsq0TtSq32erA8AL0huscLhqHJleoJJAO1h0f1EPWkz56t7RQfFBXB2fMzK3AR
a35nqQV96ja/GYOdSHxq3boLqlICy2+Y6ygLzR87dZdUReCYpRffu+zokcGFSoNIOQdOT8XVRaXm
wo7uI7RBYRDhT0yG5n//FAu3R8ocwOQ9Xyji7EE1Uigdu56w4k0/R2+sr8O1BCXN4JwxkvBIePDI
JWhDh4w63ked1BOAWZh5P5NfGc4ujlhlkl7DapZ4QIvdWSPnMHpJR7n3fshIgFqFkrXFp6JmagFS
9eI9+Iho8/MT3tOk860t0YSbJg0iR8u/n19vmXqRSqAvRliosMdCU3YxUyWLkEnOZwohbn152+jT
eBJ49oaZzEnJFuHv4mwZU17nnWRt8aDzXndbXkgmt0kv2fviU7Kn3ZhGMZqiQvsXc996SEtTH/iQ
weRLcQwAUut5hJ1DfMb5b8gxoilfsny7mlgwdiNZnxW1nsx0Kmf7JDejskkmFOw8iod4czREdURu
X3JuvLI8uLeXm2npTmbj00Mhn3wBUeCVK/MA6by90vrbZ+547+mGdj84rTlySCNOZJ8bTCQrcaLV
phGRuC1cT3AOEujEYOx2vx5HydlaHkx73SXRPMUfUPpG/CFDrnUclmizyNzdKvBK2hpJRRcEA/Xk
Vh6zrJ1edrQwFXrnXJmuXnlAHPnkOn1mvfnhiFqJrKzL8MGAFtpDfqjjyMkU28J3G/m+2X2hZBdU
/CTeSAdy7HdtZS8cS+UY8JX0zUqNp71AJi8eFGYvRqujs5k08518U8uyNTxK5eOb5mzjxV+TCDuG
CObU49Oz2CWWqM/yI0NK9CLgrxRyy80+/mWB43+ajIVzV1mxCeJ82ce0MFbBmu+Dtg2C9oj32C97
wLnXFzMlTx6DMcjlMfJK3AiZN8smMXc9CsSdvR/OmHZhfxQCOEVl8YqGwdbVmwzEJb/EtDNLiQq2
lwkZUUd1XSiWcoIg8HP1mjRPyM5nSorJuw/+ywBGTwVcsuXy0wDGA1hK8KZq7Irbg2+9tMCBdRnZ
xlW4o8bX34tQQ/L6L2NUGVjbgjsL43E2Kj2xQ+D0HxJ/tNFB+QH9PkfLqj8gRQVddzTM1kp9X28b
ThiDkwLjTLxEz5oY3W5NDMfpobZN9mt8XDHfyJSJJ9yR0vXAOIRPKAmRG7hPGmPsJu79/tB8INwT
gktfVfeUuYVlUUWEpsxHGDNkW56tMcECJ0v2B2IhJkvmkHavXcP/zzuuXev5SOYYtmUR7tsweS8S
ZMkRgkn5crXwlOoRjuj7ZnWbF/eQekAGK0XEHoff5n1qXU4GuyihtxS4SX62xWB8qQVXntYfNxWo
hkWU6xfDPmDKO6ZY6Ht74uDasqCrR+8e4aJhlsQiM4u3pVjrKAbtyijqEUPRFSc4uU1i2krJzxV7
jWj/UpFuJYKzk9DBhb2JeEPUdykwVFGTVy+is9ruMkfULEC4IBO41RoshVx2BWxBk5X9EEJn3/oI
/VkbQu/0uguvHDLQL8L9RCWdTrMzRkxfMTn+m0FZMJ7FBB6LkAlmUa9PyJFvKW0XYAdh28jgugvq
gPdNXmkEYK+KDX+d8Uw0HcpfsuKD/EatDdXaJ6to8DtDqAD2rFhgwSPip61+mBrd+smP/3aXsVnm
OtfvjRTT2/LXqshQsLn5+n8l0gP27vjfeEpLKe/dwU584PcjuDWaTj2rI1RPkcdRJRtkqEXcJjY9
m3r8mnI8Vl6AMQxcrSxYekFWKyn3UPvcAYTTbt7ACjCIwI0BXtXvJJfYldQZb7R/uymH36/D33wd
0FIHrK2FsHL+p7fPtjODWtSA7KdyEM3eiNQV26uL2GoTMzS3AWXHiRZ9imEOeL7n5HATuHemyPWl
8y5CXXyPIJFaQ96g8RbMGEK0wNaFppt7M/xbtjoOdrl0q+KT5BIq+uoLWotND6UHRj7PVDAjK/D5
D5k9C8i0EyiBnnIzxBFVV5+d+vStzCOFMbGqPbkf6at15fxGh6kGX8i2zI9FRKk+GvFT3vmCCtEg
VZKLuxgqsRDmRJZuSjZ9Uieaa5hPlxbTL31JPu1nJT/jYL90IVlu6Uz0hHnLBXb/xVS7t0Id95/G
d1/t9TP21Frhh7tv0p2uSFi5OJF1ETgaDAs7B3cai+EebG/Nt0t7hS9EjiPadHoRsFaeouXgkjaf
Nbh2NcBBN9eamPEKKC/tkl3jc0rfrUNcSdofENEvI1049tUTUQkRMZ60RTKrLzuOpNReerLNhpok
ds8RMd6AMk5CQoYz9tRs+hnddFlmCE0GiKE4wADipTUCUfDZrMC9YsB18pkzSheWxXSvK+tEeieg
VBhX9rcgL0kYdgVv0lz8wil8E4Xbj3WlCP73nmK8fVeiAGvjqFSRqxErIFEuC7HTbcHMbdpSpq9M
pZYHZLJ+tPyzTrSwCBmd/ykx9lMIa7PkS1OMduCtXcokK6kp44PfPlVPUHuul//k3A4fpxBu9ztP
nj/TU3kNfeXqvYpJs/sQvc+jvD4EihllCgpAybRfk77/TQiCuzp6e/9A18YtCAXtg+ezu4mg7LoW
KhIjEfRWkAIaIcKts3+zLz6uOozdckzrjeTItLnp0DM9vLCzM3lSPo5CXOr6v96zJDbcDqzVYYP9
G3Pg7T32Ksed18INt5dWJ6fR4ruSOxQzHKdwUp/Wy6k30e16c/qL9IfGa1Vd6tdO8NeFms6QOZn8
WyCkkFbNblYhs38dYboBwgsjNmJYv6BEmRQZjQYrUAtUH90Fr3V5YJp9HOqcPRC8AXsKb3cg3FXc
meTBXy0O2NZl8XUzeGq7DscWfQNoz5jUCq8Id+/6kIwsWG5GawGTAjGAONSs9P6kuhbgizCSFKcM
4nk/7G/dsouFmN6tKfb0BsKZpDRT8flQL+WxZbxmaLORXnkYVvUztdMigLNVUX2ONdlslLSTBepA
2dDNkHt1m784ka0SwK0kZZKv8ReS+P1ZEsFd45CP/gvc2ztsqxQDSgAB5R4Fs6z5A3wgqhQHSAya
R8J266iYkShWWlLqM+EFDflcsjt50XrF9lvRvhViVw7FPaeKE2pozEzjQ4EV6gaJLWgvjJamBae7
CRaYtF9iZAOhmbvBYv6zppSfe1E5xH2xz0FmaIl0KvaQl2Ne43DZuNQWsIq5VcyHWaenG/t6ySly
2jfDqAjlm01pWO6bLliO/oWqbvjjcpFXHW/0Ld3ndgw1TMp4R9v3T9PMcJqcz3B/11/rwsYRpEcH
ZLgpvUi0ZJ05u98w1CEvjEL5wZPWjj+GIkNT6bO6JXJ1qyIip+9LhZyIah5+9ShKB7oiPmpTeh/P
Lv+6FOIbiJTTarj6XZMOj0b4TBvx2538QsX6FGY+IE8qJrjCz+0Ps6xOKXf8sRzIIZVaL9pjHbKi
jUQeKxdu1CCcO58ynBQ3Y1h7MA52b+qxWeQQmB9OAhhrzHFJ81IlBZsdyvtXgSCe9o69aRW/EKpp
1HE/JcLWv4+xdIIVnZFMGxlzv942Krrb/dHcgvKsicXWTrHHo7EciQ8D+bK/F+R6KERx+hb9eQ9c
oRRRxwtFj0Tixe033ZSUfoO0ybQIowhhPc86WZJJ+2pGj7vuPevhAwek/9awqonm4PnbN/PA0ixc
kl6b5gZuNwii4c3NUbS55cy3CAFE7YwmJEj8cm9um3pM5yqQ0TPSvNme53MnuJ5KITPI4kROB878
4p7qwJlZj88uiViDbJKfsXTMr1jCBIr0O7HIHQoEZ3Hz/YkQZVrpgkgxmb6BUTGa34rTK0uYrwOu
DPCoJ+I3jUHTftSqqMZP31Rg9w7PYjmNORw7dBLRKfsyTPF8O22shVon0ArJdBw/lpDucV0Y6yDT
WWyujVTlqA4/l+XKK8aBSE6q4BaHo/A6Wy4tjtWuwDRcNfVuGzXTVQas0BzpxOk2VhRLeO4nsP3M
F3FM+j27uvL78GVo+kMuy1zWOM1V3zXwQ2j8Y8HBFGf57jAdPRXERF8okZtr0R2wN1KEyUO38pIy
hqKiMnt84EvLpjgWzpD+1RFRPARH7+FNgk29MYfrQUAG3RDnANPXuS1An8OoJcp/nB/7sAHT/+W+
A2XFcQITrB4dME6AJCgjnxVRMJBDt/6wZLCcUffHNfwcPMe/ynaDKw8TRejZ0Epf4/VTmaQ5ZGRT
rK2jhSyhcSwRxD6QE8un6A/wsPgeTNFJRuZW3kL0Wu3khgk5mcby+2EOULAMieqHvnR+i1Pa7qQf
YdSU/6M9fNfUFIggMIPFmwisFYBn6Q+h7cKdWCXtPffzZp/+anKbkkTAxMczMfki/rOmsSIGx4ns
shUzu61DV9c3tseUt4pJs+OMwGvBdggjjr7N2goPC9g+eqsDh6KlMoHsmGIO/xeoHZfs7YxhS4ye
Fs0p6aiV1fS6F7wHJUrJlJCbFDwA0ToJ9hbBanOgrxgjPeAkchQWlEswh5oTS2JPgm6JjqHPQqvy
xaeCUeyqCw9V4U/a9brWz3gS2iHZdZevk3WyZD6L4ee8WKmn8TC1Nci70+k2yOr0oLPzTj0PZNZm
Vvl0ezt/pVe0yyxQTr31LNrdliUnOcUuwXI4/kE93QtBnhgfEI1JR/h1gsPJ/6+qN2ikmNnOHZA0
4Leza4xsA7YzmjQwlchAKHUvDRnQ06f4TpxH7mCaPWf10xnbGZwdFwsntT7ajrT6rF9DphbcCxPj
v1A/YHnJiW7/B+aN+W8BDM1gUIG1rFbRWK8XlJcrb304LrgHVjZrcHCcKWMqnaciZdAyNvptr9Ju
BTF6iC8KazanR9WSsNUPF6o+TA2Pf2pu+y2fG6tc7nHhMJXVvvQhMR58iHbMbt8d4GhxzrDnm7Hw
b+Li6HJZvtzmyMw9IMWVojU6BjIXD6ARfIGQR9eXHAzaBWIEcBEbMyIh4vR+Mn6YMWhfuZTcCTg/
SIzl8pd/1vmrWU9jqAk/tVfDGEx1/KJnnrD5ka8aTaG+TfVsLOVDT704nfRZo+7dhl/GU5hVxUUn
JlgTWnM9E8H6asrBdK+7BINrFBxaUaNlvGKaWCD+DmQb7R9z91pdvxQsowY293ZLWmJWFc7foaFZ
X+F6dZ3H4UJlV90djArTczF5bMXuBfHWqGkrjhrntaU6sbzuAHw8wtalVtJGpi8VDO6++AvKR4fB
O+55+RPeoa3WTZiI2AzwmGrDBJmmBa2f41Gu5JVxgs2dA9gLG8+B7F1aGBU0W/jqESjw3Ltyzows
LbuOSNzBp1u5N+n+3CCfDRGE8ao1+5Tt2O7DqwhW2eyE83WQobGRbbHx495E6sFINsQHNlqP5mOU
Qy0gyZ7NBtmpn++nlN4iFyiNm3t2OQIPXPdWHkRvlfbsRa3uRqrfQVe8v0hvA+UsajGQgKKkXUvG
CmOlC4TZM5WIKKqXzDwtKv7aB3YdIhEY8o9sdAROLKqXO+30RIQ0nSmPejIbi439SlGCxImcRUW4
wH2cfYG8djH4r16Y8Z/+n6VTPzH0DtZqD+Y3Sbn7RK/w1Aw325UwGCK1gRQkU/3xZNRbuGJtgw/a
s6rnAThk++kSuaLMIkCldxtqIXWAJ4Ba6lPUWaEGmw68b6+D3yRm6JS3kLpEKmZJGfrZR7ecO29s
ZfcrlDti5W5LanSsFuCTzJ3aZiWeeBObUXOVEgJS2/f5SqcxOXKBACHb+ix89C1dXY/ELvFo/TiC
7qvZ4cXRHSxDXbQe6RtNniMLfupvuoHnAH2lM6/e6fEpzOZmii+B9YBaBoLCsB1Qbcl2ovP4AlBM
czaqaCg56kZlwiHuuyHoGPEZlkyf6D0CaMaOHmLgBNEeUOwIMuayIQwsubRCjGKnIcQ+729ODcqg
kHe53GMUIcS49mxzl8x1Oak4QHthz3OmF9f3hsrFLx37bpXfkU8aUCb6/h5E6LRR5P1KOLGIRHqN
gBFE6Oe0XFthrR6jyS2fKDZGJp8yqksaeHhkSLcTkp8KFfKcxror6dmWhcz54vr6/ko78/MBNbE0
1G8g5Ssn2QfrkKNdPkL1hcWukxPb27p2uBRQtTs0IGx+yPQjrUt1ngpTRx8h7VfhEDv3EUSu8JEM
NfwTA4mDar5KZWUmfS/RI6FmST0BMuO5zkL8MS0DDu1H6bkm34lQ+cakb4rdFPbE4m+3HWx22diD
sLgtmpYvfReLHoWS0HpjXykUSZl7Z2b0cUDC8CMxq2C15DGbh7fm+v5km2qwefvGbzbNaCmnXXAc
Ws5padKBFbZB1j2E53E08n+e5NI+qSgHAeuwGYU2P/A+7sUVC5ZqqCSdE25jmhEuKObpEbpS2alq
dNTU4Kx4ijAM9TuMVJxxbP+ReCsT1ca34VwWwuJX0TCsFgW0SaBX0YxgTEeajYyiMdpk6LrjXxzT
JiX9Hzeko5kDQkjlr+gS5wjgGfHehWvj3Xho5YeOCB59LzD5eNbM3/YQxrodoHdUAbjKK/zFYrs/
IVFhfpCitMLlLbbEm873EAPErRbytkcy2ub6I7amOrLpGQLTaKqu5g9izm81qkoUsyNWX6vK5acC
X0c5qEWAH5R6v5F5SdYidg4tL3FR1jp/IQwrq6c2J/9Nllyi3VcvXFCuMfikN4dXcP11rzgkftw6
nTxy0l0gfmm4dFJ2RlFmRwwsc7cx7WcZTuDxtmw4YnwNkG6MrsPHtfWg6M/SZSIFVN1nR74CthP6
PpaXosqYo+qv1GCP6v8dbKgzdorHTfUhI0mwiUJz2//qBCAogsHaLR3LnwBInt0Oz9OQXXJY24qO
tdzdr4klOnVbK4cnudL0W2rY2tOo5123uMbOyrJs9NeZk6FlWrKJ1cB2bIzIrBHhXRprCbZqqnuj
dYvgnt89eIp4IxOWXTzz1DA00CA/jXYKXDMHxXCY7x0Lylc4yeusscI4b4NDWS/E9sYYBWt0zSyi
48lRH838SeYPk/u0klA4JN7E1JYf9OJOxH/JG+gDpJh3GnqeGFaxEdPve16BG01sG5yJAA5al2aF
B/IWODv3qOQEMKnQhDv06NTdjDIga4Q9ku+i3G14eYFBF3JXJYKoWbF5MzdYc0I0/NVSrePI4uxR
ntUhEodEo7Rv3n+9oEsM/yhyubrl9Y3IAr/D811nTdq0MES11seAfFP34ZZbaYQuIKX8CFw96bJO
4Rx8SQ1FvrPvSBZgRrBZ2SLVFPUrl7dwrNB38Em8hAkOQbdZaHlHBwEbMK+v8z/uSfwyGE07dns0
1bKRUOO1Y7F9b/cUTChkLLXZ7jJrNW9Mbbts0z0Y3MlR+ApP1L9kRwdtYrPz3AQ6BmD78cRX77Ss
KE05g1F4kHRgP8xC/IRdAvT4NW32q4xk35ge5Q/vC6594wok4Xfu+u/z7wLAvZh0Dn6mrYjFGxbI
pLD6/u03wT2nuhuo/3k1b7/uDbqHDZBt+w0J0LlKk/dyukTQuihoWqRaMr+lEwQUsNHs7th/+LW5
u5M9FNeCiCPFRxGl+iz0GpNd1f1xyNX6iGQRrQ0YtOYCIGc+ojd6nPRiZBXVJc+DOpSymGjg84XO
ook+QQpJoemj+KS0Thuodno/3QhDucI38RWVgS4eJO8QzkHiWnaUwxqcu3ixMV7EcsIDTjLREmop
FvoxnCKqlPHfV+ZXt6ZsWU3qv2p7SEsAdARSpVf+BUpF+trCLMRtQNl2VuFmfhBJ+TlD7LNr7zA5
BQyfyhI4URl+fu8XH3cNEqSOsEVwqpCzVbqsT75YoNdDUF9AbtTkHUavr3Lc/QGLpc0cctveVTE5
8exxZcOFHao5xRtmGnNV1XmtbrU26b/m+sZSV+biiW2aEzChIa7K5BZ4ewbi8ox2mrEc7N7HP5Dz
tNIuH2IZmul9Jw6rfR9KeP2Tk2QcmNbrwzecgeW9AE184CiPhPUmyth/Iy8/14+KzgrK10cRnRh3
R82ghRvuStJ+xgbzq0qrNL05E943oj2ouhR2crhsCx1Es6Xfl2CQAVzjwfMYx2IFYoX2jDOwmcly
yX+nO7k1FKTj+fGQEY0q4+XLnUF04iHuG1lQV8QRsQoNSD+u13ccMGCNL9fHVc0FbQ252N7aokQo
Lg7LrQPAf6cBHrYmokMAeh/y8xXaOwqo5grIZKL6SEqhSGWt/jeQqLvBE1I22CbeaENvHbo5Boid
xDqMfeQZsNi/hLz9FJUiwbkyBUYKR2KcNiDj96DVn4rfYXIbSgnZ1hrJ7gLq6z7ZWBvS/a0XMeJC
lEooHcpyw5EeEF09beg0EfT2qgtBn3DsWP63jl3fT0q5MAunHTLx14U4My2B09Skg1fiMloojKFB
eTyrW6h64AcsPQNch1aMznDCmRT9W6KfGA9poISC6vDUZzZSIIBtG1kLyAMnBX3UBB6AAwizuZuK
YIq9rWhjL++AAd18g1fAM6PA4TmF0NXlRtR3i6Zqd9OLQ3I5pEowB6uYuVRm1HBopW9+eM6TDa+x
P70Jx9F7pzeYjTOeEDMyBtezwNLVliuvyKRYcwyfvNKcD6NHDxUVfaBQtDD8wnzfF5w2EsZXERvr
UDArSWcaEYKDCTSSDgCTF9Fc4ygLSbRd+z+9UAhsV9ECsrwGQICLtmFWnCyuK7o5RmMnGNjcVMgP
Co50jMphAJWKTA7+/8hzqesEbshwYSOZCnpSyHAv3ivuVKLxCmAKprtstPp45PO2URqHJZZhb96g
r2dxsF6eWi4RudnUHGSnnB0SwNiLZAXQM3+efthKwg6GjNUZEoxVi5O8iJpG/zgPC1Vvxk2xenu8
cbdPYlf4G6Bgteem2lTPom1s88X1Hn/PgvWS6bVYgvVPG7GODZf9aXxStkk/sLb1zDTw1tu8EyvJ
qwYBkCZ7DqmY+lBAA2mJPJgiAttP2ahTfWe8YElUheNt2EQyiUc6td46nr21tON+TxvudH15pOfw
roEZLhdtGq2rjDyIddnq6gdWGuSCutWNLqnfhgs8l7Fkb8czaXM0lEP9VIWNXR/UzzYIlfR0Yp4q
ENNGgurDCp2e/GNrdA5GDlXcO9IUD7z9nMWoEZUKYeU6Yl4kakQcqWpB1mhqwzIdPRvwkJKB4CJJ
7NJvVdwzwrmZZHev6Nd3m6tKScFWQgsr4sohvShsL4pzYfetGuEnpv2EfabhH5FsOHzuIBKkDCrP
I7yOfh9yyT9zrTK+3zlhxMpcibSz/rPGZvxiaZBvouZZgj3L8AmQx3zcxESdNfs4y+Z8RXAIkdAj
AJKxkUcinH7p5/Oi+tAEvhGXFxppus9DHAJqEPmJZOTRBURRdSCIN7uGkQQFMpre7wXdOEANNZvl
dTSVr1/BDxe98hqzMl/qTt50xDv7b6Oo6Ipou+PfmGWa9dLMmhqV/Dz86FPFAMToPDXuAhozO9Cb
36EI6WpwQR9PSxvCx4IDxTDtnydPzq/ttiRI0Mx5lKDoklPE0+wrmHJPk14NlsbjOAyhDIqZ+4X8
A4fQtpX6iVgvXCii1AaatJXDGwoZssfMwV/PE8k83q3FUcSKyWlw6EyMO2hsuqeYo6nNlBUUB1X2
hxHsiVQBb/OEtegA/jzI2NPwW1z1LvsRRl0TTYt5Dy9vEuNRT1FC0QRZOtmgZ46ymhsYO3kgW1pU
zKb5hyk8Bg0jcUHIoQgntYH4CsskQflibgZ5Ii4VYbp8v479qEP3czGedglZa+CKEJeDhT7iZodv
r2tk/55tz7GiU2q8Q1xKpAYgODbEwtuV9jyDNhlDQnwN9tIp0oW1ToGhyAdaEBhsB6GNo2Bgq53R
ze1UYaC+DB1r6F3aTP0IKWPIsY3vyri11+JOtqJ3fwJp88CZqygTPWjph1pbPbEdD/MxTjKcVI8Z
puf5kFmMh1lwvaREkyv5/sqKeuhajtjPTKLBLBSEyFZ4Qyn9HzvmQ8jFW/KTaRPeqwvC2nNX5gj6
3rayBBKqRIRVqNVirKGpXLPpERycbU5lAGC+Zdn52HszfJ3kxmlPsPIGJSZNR9iTMqpfqgFUkI0F
aAt3VOXEkO9E1yqkbfoVCAcPWTg2S4B/pxWHFUowBpbgc2TTzU/Yp8u7VVDoNv1eK5uUA3FV+qya
hTtm04bKoITnnh7k1NsKGKCNc9b+7RGEJLz9DsZORBJaTLlnLRgTQLlVLVTLSBrUDLu9+3CGkXYF
EN3vE3COn6PF70N5KBAWi6tq++mDEjuFWIe43Jlo7tNQS2RWK7GblQVYyyDPLbtA5eSzH2bwNyWm
zEzJeeHq4QjT/6rJ9W7BwbTg/x0q48UxQU7k0odCmYOL9NkVhmoL050ck7H9RSp5rSBXgMQ2PCQS
uw+7zxrrdd8FqeowMSzB35L025YnY6mhTAybJq+idNYIpJivreghREQcPFR4D11J2SXcK+GGng3K
HujjlxA5OllLHG6QyC1GyymbmESe6cLPggqxR+Y7kMnIF1acIYMISeziHh8PR2enoBIT0SvLXwvt
OINLZxCGU8jESqmiCrwt90qnmlqDmZDQNIkUPgYVog4ceurVKKlScGiQil1VnyU83XcAQI5+ER7j
3VSxMwJ3X+OKOMlqPRuP91FtCVlPLpMaL2oSH8q4eYSvDBE/joc9HA0Te1/q7FIoLJ9x83QDUmM4
ndfHBu4jnWp86Gc+nG3J4IBywdgHjX0oeW6Ppzd+IemfM3889ss2BC32Vo5pNSr5PrB2huz5PCcZ
h6KtUTwuWSGTnZ8TFMPw22jQgAVFePWdlET0wKuAbj/w2lrDczGL8P5BAfJd6eiRTWOC+dVGBWzB
xOer8DvislZIyBAOMVgBoaBuRwRH1Fs4Z0r9+QuTXQYFO9wBmqYvQQqlz1oAB+4qpVGxCVFKkVDA
UyTt2JRnHJlqZzaF2S4nD3QAl4v6vPwvDrVOAl6WOZdUIOtKL0Ebo9eE2Tt8WyIvUDxdYa6VoQeJ
SyBoEGh/g7yjxXtwM5teooMEqThcdV7/56BRXS9PQYV2t5K84bq7bYvqka9Aoulo4aRQy17aq1RA
NPUJsEBMMtkYu0iLABW7npECN4/2HnrNDj0p4cESNXV8hd00yloSpGTmYqBJQnIlJ6QtO6bGiZiM
N5ApD2js2J3YSCIhHFdqYWud7hDyMQXdh1Aee3PXr1PyJjxpPOaPSiCTDMHEZ4yme/yyezboOcnp
ELP3ysf3ie0oQyLELjK2y/Gca+9UTLusSx4g1pAKjRl1UK6UqBQpbmG2XEFcVwlX10u3AtXzBiis
t6pzdOOz3SbSBeNeE1SpCO2mvf4ntLsEbYPJBGjpzBlDWMKOnjG+B57NEOyk8pqA6G/HlJ63UO1L
JcJpN4H3FdTG37MSLRunFjNlA5DNp6Bej1Q4yUoAljOzwe7Dao/vkyV2XVtCtRMOrlG/yFovg1YT
cyifCvwFoD8PSN8CCeDz/Hmby3G8+KZ2NjESRMZY3l13lLtoF47VK9jXUc6T5XekeP/TqFkBOa7/
YpyPyHDB+orAkdFUMiuNd9IXMwvG0DMCTuIZkClsmEfc7Z+9jYJ9qTZZqGUOilKg7u6SFRS1o7jQ
872c9WZ4QCsW1lXYMCCgst8dBVH1cTsFN1wwWDRoYEUPFNaF+AbqoWiQIz/S/tNiPnqtD5B7i/Ci
Ueb1BhGPmukQl9sfpfpCxIUlhdkbl1WgAO88b7JhVY+BLH88+TokGJYJHha4/iqRs0N5ZJ+1VDf+
LS64CUeZlsu2pctiM6+1V3u1rn+Upb6pKtuJXlomy6bwDGLvsfuGm/qYmKO5xI35r+AIOJE8wIj7
zoRrSwq2n0qFRSNI37tsh3zLP6u+9RNHC+lnx2X09Rh8XfBDbw/qaFRb2MjWmYFlFHbavFxR9Gxw
yGzmsacjiZkx4IHa2LZC4nTANtgfO/GoMsPZJiZfR5AU5DhMI8Nv9JVeR/tVnfPTM+y8gIS03mOo
G8LzesnCCwPPFUqeFmBR+9NkL25KO7IqB3sorFba2OydB5Cr3MNZ02lMPM2D99c0Q61M/JTPh/q/
ATS0J8tjZai0zDIC5oEbTHb8osCrlxEp2O283Tq9uD571QHrMDS1lA4LlRSRQtv/eDW/XkiGrHKQ
ttNMVyA/qRMLPfeZcIuXTvAthhkkPRi0hv4+6HEHg/AoD8Rd1eIPN1FtgaP64aXrTy9ffEqrcPHw
z/SOwGaAriC6CWYAaKbeE64dEAcF9G+KVfBDtQMwW5QhQFLy8U43KNefdLTLdtOfdjCyWIdFvpd0
zyUJ84j5Tfg22RKB7OuGb+SIeDK+E2jhLq+bD2Ch5rOwuOFF0vFi49VJKZykk27gkms6x+LqcLQz
KopvmDmSgoi2aZWyoqrKRdkE1A2rQcfYoq099qOTDOx4U8pkfXoH5MrAHhTLHQJ1LeBe/HQ6KsZr
L7BJ8fkB7ufOBXrwbJY3aWPkVD6feGnwFSsZt57dinkuK9gsc3AIKAAT9Ogw6kFHsAIjKBIsDGfb
2jg3JAou0V/3zQjdlxs0LAPkN34Cu+HSOAZg/gunGOsaIm3xuoRtLJ8ItPeBRFxfavNUyPwOyXZa
Q2bdvqZ7Yr1SizWWHUgHrGpFlDeY5Ewx9tBldL6Gvuq02QDTNve/xMQ7a5USgtVtcWsjsy2aCaVG
mkrqshpMWUZ2+0fkts7haECHbDwzLPoaD1sRNJp/d+22YwEv9iRarZDoZaT9n+OOUyb2Nvt0Ze1D
yMygyBY4z09i5Wsv5VP2fObylmfEDkBfYFdVx2w/W+PpcMzqAdEmkYi9MW6X8hmzCjEVDUD/vHNR
tggDZBjclU+pZ3iArei0UtZop1PYncyUT3tUnaeCFUibHyj7C/JnCuzqdfKuLCARwr19jvJSJ4Tf
MvZnGTdJF17lSSs4eOFzmV+S58eBwV0ftz2klZf4kZdQSVGuLh+rdjBkONmg1j3vQJjSMYOUD/Ld
s/0mIFzQUguhWBQYysIdtFILo1r3s9jBWnIGaCXgayaGnwle72IFSnEWcKb05aOVpOTvGGeruoMJ
wc6xbHb7YvtNdTPouionezXWuvsGgsbcNr5HfIqLv6dQHOnHNRXZGV9Kn2nuRH5t7lXntXF0yMEc
RYPzXnkZENxxRs5b1GAzhRjUG4FtC+yNzV3Y1NbyWGLiffwAtjX9rb1GYUSuV96xE1X3AiBGJMM7
rgv49HZPz8Wzxb+jgzQZVkYyUOuZ7ggfFNDFSfAH+w6dG51dVnnP2dGJTUAAgQv82iLcTI8pe41D
FnNFNKP/YgXeQ6pwy5joCPMEBRP9Avb5rCR2JBxpBjoX4fwG3sDgcsHIh83QOE/y/FqRPtJPTVzZ
NrXhe/O849DyxFkZtJjP922F1YAH5YgBBut0OQAjCIG5NmRmR58Q22+u12gbJFhOYvFRt2KpC5ou
ffWsuKxNGv1+Y9sOVWOchEDhXFdDyTsMZ+TGSlo2zxk/vQg7a3v0vROOL35hBpHd/Trqr39EyKRd
dyd8+TTHnF40SyK7sVI8rBW7x2Reh2pzB6fT5dJmp6/TzhKhJ4gnKStwsGmmu7fh+7lqLAB5zWOy
zTUOT85hKxfxQfvrCMKf4toCzasEKoL3dbZ3YpeSEWsJw6TSOxeg8cAXK9jOrLFlh6pjWGgmuzPd
kzcYKuW4mcPz2vKSTY5n+HgvODJhHkupsim0ZRnq5JxuqoCmDopPB8Ydn4ySqPj7qc3LWZThViGe
6rsCbCxkgn9SvXgQkcQ8lE7OYfydgMGCJQvj/VYYJFQEvFBUbl7Xa1hyZzDzPWSF39n1uxj6c1iq
F9x3NeHHuu2VKGkfsbHbVtGWAXY1/+kMbdLl51Iggtws924BgOkQ/r6LB+YnmAIrK/o0T3g4NxTB
8VBwL+AV27XrPvVrtBJgWL7gSgHhVU9HK4eAjUP5f3YeL56T/Fm1wGOQk5KhoXRd3K7bVP0ZD+Rq
TxHiNGeLqmUUcUq3iQgW38XYou9fyov7xUhURBHWIkZiMLEQu7jobVFsCp5fxqTq43tcBHx/3nqI
aeeXg98QDVS/iV0AW5/MRC8yxvwlfRRTN40rmxP5fXKYjCcaCJuCSVWXpoG5rBz8PHhuJvo41LpC
AJwK2PjiR8MqubU8W3PrO6LD7o8lY0KBQERjS0NHmIno6cXBlANpweB3oHbN2nsCtrDyHkiStmdY
qYHFyPIWcFJUeNOJosFw0ruxfhMgaGhiyzqwrk0q5m5ItraPGGtPPwwFy6eRlstQzJxLEyPPwzJv
Dx38qw8iHqsEJ/IOp2gTiy+7OloJxolwZBJbVj1s9v2bSxHenf4dt9Go2YRbf464jPE/IeuVXJ6X
aV73deTIbREQmjDGI25CI82XQH4JTLvmqSULmCLsF/EQapE2y6NgpvH+0qcz8GXew0v0FFf4VXsY
9Th0P3/1nTO6X1/xVRjjwYi0N23NAhDbuPqGqzfgkPt4KB+4kZTlTRePZDvvbSMoip8SQoHhNuoE
jSMgn7rBoNzvMOwFcefprvyJTILwgkMc/nKReQyEn2QqqJJYmaMB7RxdhNYvDBkBKNCJkGBZitki
v8W8w2wvrL/0BM5QF34YK0oJgKh6EV9cMsJKIKW/mKg6dMFbX3Y0AtW81zgu48HN9xNP8j0d896i
aSNEbZr0nwDyw4MKw8erfjRU23cLrijoG2hVM1jfFBgT6ZAI1ORS/JO4gHhP6AltxQZvnTy8Tzv6
4clTAfNlSEiFhaGxRj4YixJCQdK+IDWCwymLs4ENZyUIBZNb/xmZqjY1zJij/KucbP753XlTCYlf
xU1pZ+Nzob9WZE+BIq5mTOJSwsDAQOvf0m2TcpDUpACvDdO3Kgd0zdJSFq+sPHFnXDPzCsGsuVEC
F6ueQPMDa4ucOXrY7IuBOUnkCgFPLE12h3Rg/lP4SoneqUuoPIGWoTz5VfEzb+uRrMScD1QzrtV5
QWocDHtWbg6FmSzXb5JX/Gr+3xB84fhxWkZQOemWwBNjKwpYbTy3eeAU+ByF7G6rmtuyuPhcapAM
z2QkBrlrSIeDYa4RI7yyOxgvxsnq3MMVGlLAkAEQBhKQP3mPjDvtu9X4Y5bTF0RDRClyfIodsd/T
UyWdABGsDclnfLgHZFk2peLo97w9a9w9itWHMnWPsg2lXTB8i9Hm+AmaXdAlLvM8cyA3uwLoSVYN
JTRIUR+HMLGUals4YIHWl1Civu/OWSOwX3QxDBf6xX8LZ+sPA7NJVydiGNT+1ku2DkoiU2l1pASt
N5UwiwP+BNgWAvxdjokPXQCD411CXyzqcmXqiGDUK3hhJ5Fx7+aODfUzs8GGD89LtsD4KxXn1zQf
Z5Kj7eFJ6lSp9u9zUAOh3rs2DAUrEzKv0HkrDXl1Rbc4KMpMel50dndFieX9oA1v4XYZiNNci0sx
xFG795vLmUlx6NrZGEuMdy3Ba1GOCb9/oORzsl/gnKAUxjTJLRO+l1JaqD6pCSDsFuyLPq7WTQ8k
CyhZwbHqLTavmpxwZ51hnLh7aK5LPia5RYERXS+K2Lvrz928p2SSTJ96Ct0LZGm2hiszBX0re+/U
0+MSn3tjg5dTbY5MSnNlfTsgOtk09ckU3ywfvg2Aq4DiWruI+qbztpX0KjIXnJ2pJ/pDP4PmHRfo
MMkISw/rTwYP38rOHcldpsT9V1uBOgTVj/K4VSLaWmpntuYwDkkfLOgwku+ZIVzYBlRjctt2ZW/E
gJyscUiouCylSKroA65JL0OFaNgY06sslYSaezZUe17lqEEasCDT3a8UZ08eQ34GTYTkIg+mnPMt
uybN2/B678f2wyD/JR7LDleoBEh7EMVHTKDScFiaDrQbZUwGsccQtBiT0pjrctl/kasIfbl6LBi4
8+YCoOfDmCMVFnjd51i478D8gYgOsp5d3a8AsdhkXWjwKf98wYzIVUJj5zlm/7VfJfo5BFVou//j
7Ycc5qTCVZFkPD3pK9RBpCFwo0mnvsjc+8PjsT2jgzPlZngkQVO4JbOBTFDtavWmT1u2LCjzOrjp
Zw/rlV2QuQ0YeJWdanCOA/QXVmMsGWNQsfhcZyGeLaS3+qojvv54JTvVtWDGgMjInPQQa401sO4A
d1ayNsYvcoRqq//w6sxqtL905H4Zzfw4JE0ra+70FxyyXJ7HMnkZmA9KeXqFbmPI0dQbZ/YuLocq
vNuTStqo2uL2cGU8du3YV6PrzgiM5DmBQUVTfq7ywmU1G9wDBGgObRPkrw8Gy/jnbU60U5atjvtC
LdO3pd0YkKn+20RI220Z08bgr4n5szHABVkO/M0nnfe+k/8KkZQkaa28bGabg5VXgwSSN5ghIVWb
M6W0u/Bllfom/1Xvu7XgyYSmqUqPVw09PJMljCCBrS3nighpt4rFTIxhmv17OkvpeeDFtkxavsUH
Rly9encrW6ixknscVEULbL4XylhpUECwjoYC8PbeuppXvwl+U3CKsFeXhBU8D4gMf+Bzz1aOxb2f
T84TGz+MKC7/7EJrUSkIeHN+ix2cXY2eOUA6MZSYBfo4xomoTwOS6sdIvru2QDrZurv9rf5bLALt
r8gZ1Gf3vqQ7IxqFahXzy6ZPJFDxWyeNHKWy+pDWb4aOhHMNCQhbGLQva7wW1ClYPtkMiES+trWP
7k1R5inywOrpV6NQPBmLPnii61rQT53g61A+a28cqt/6RyFJsSw/iu/EZw4j0nLQAG/oHoyx7ax6
bDOESDxWffdP4hP4HuaG0u1KCIgU15ECVCl5NrGfHdi/RSGmD0nk/Z5DNg7Ih5kUljyfWwn4cVd/
kEJUj9c59LPDT7QVgtaIb87bp8k1F1otzBG8AuUVD+VYSHB4vfUmxR1EWxHUFNIm0E3NDX47Diae
hLBtkLAz1haqZqbqul5sBMLtBdIte6U4N+25MOj86T7dfGw5L7uosbNTmo1psCuTYGIVx/ZKE6W2
7nZdBwKJ1iTb9GF8ugxjHDqkPpu6TBE/wCYC1HX0brZL+zuDjpjHrYcbPgM+0QPNJwFKS2LZIVl3
kJvmAxbft+4SUQTZ/vC4PXHlS0V0Z36KTg/S7Go2hYiDK5vfVdn+L4DCigU2j0UQQzEG9sJbwpoj
N2h/qF9yMWFwRX1Yiyjb62+KGYHl12xsdBDHzJoVmPLBCZkTffUtpVbLY+DOCauwT3iiYnDnWmSx
syFygYZ48ACQEZ1dy4JStkKRwH4QssLWJmRyAvo0n1lLJ5jeyvLKpBr5CIVCC7Lp6xE9HtqY8WjQ
iKBl1qmO7dDlggzBj/HjIvZEhKfCXDCAnnwEc3NO/6mwiWk/GtZdVgqtP4ZfZ3rvuGa7XW1eFiaF
vopbpr8LMgKIqhiSWyqMpeOgfmIL1N0W+agA+E2wAEICXF0kebI/fseWYMIk4FtMfqF51tnBe2ys
B9xRK2VQq9q1gW5kYpqtMxjFes+KusBRnPoQbUtXzGGgHvPVXFDXDbiN9Qerbu2dctNqqQSKsXu/
05K447ObjydDG30I6Ycm10H+xxjt0FVwie+Rbb3pYxV6tBsJ8Vm5sy68Sn+1eZGVRxeKElN6TFo7
LlMofU3pzGj8R/mCHY8qjKhWHYpFNlmIFeefLWUUTebujuz+a3KP48o6lYZ6ShT0jUtqDMYLO8MQ
PWmqpzVx9gdb9RwmpKa8Ywe5zp6xjt5lVvZtAeVOr+1HkFmA5Ke3LX9XcCJTlN2yowzjWVk0TLpC
h0EkHD92ORU/I8ciNvp/U+TA1LGjC0mOxebZ8azLfUJXFSTWqlCz8EcEyTuZYogjN2Ym8OF+iIXg
CAVwcaRsDuu4maG9qRYC6DOnL70rOcwpab/o/8/DbWjMUGz7MXdIN/TeU6bochWv5ydcRxxnKoZm
am56lfvqsBCX5Na+UwUyRtIApG9cxOpHNjPAS35vN7GBMLeRl6+p5F4joUlTmm+7vWeudb2V1mmU
+dFVAC6KJpuXFiAxnaOqrADLdzRrWARySATjcIW20kRv0UoZAcQpMw2x2d0rzPsmGFfXkx9hLqFE
J9z/gXJKv0z7g9XIwmRPdlE8eLbDBn/swrbPQI46yJ0yOlVfoRiq/O4S0jpOU9LMoGPNTgDm/YWr
W0t6fjFpGhioa6UEpmZilpFZLTLvmkOCd8eGTATWIvLUZBoyaczrJx+fMFnccjvPyu1RetiDXTT0
nHhp4E9xwHrEypkx0Z0oz78aDwXex4NXFpyLN2bxd2J53ZhV3Ha1IKAMmKYMWDIu4lfAEn8z5QtO
Zn33xX2dAJLfJdDR0OlgTbLg2uJWzE3xn0JDmWHg3CdBRc8ygYnCzR51Dypq0U8yMfR1zbQ6R9HH
dtSfbs7Mpaq0obG8Nar1uFL8TlIsVnDxKlM9PXTA0SVwBbj3wjplA7tKXBr4bf0UcEI7nROrhoWN
pCVqHG5s+nMelqNTBdFVft9XKD1NHErSYUIzzQByqxnRe38gacnOA1M2CD62ffCC2EUh0k65hODu
tGyFsaKTiz2sTFtYm8jah9rocVqp0547fsogacxRnrHTDKuKEWtmpjDQ3QlqET8w4RawaSe9QZQr
r2XqlNrdRC15TdNZPpvifI74NdBTg3OFEFs8Pl7F+rh47OiKXfiuFO205EEc0qsx6FpJ0mY3z9AX
/9TriG9QfB6uw21xpcp8hwZDc0C3eL4VRExxjvJmzF3WxiQsXu8PujYoYkDYI+1EvejfstLai06j
CedArWUIQmYSUF90TwQNrECGMq+qMr7Ou+aYWhaF5r4kaHJPIOc9lVrqpY/5MGIg2VTwQT8x92d7
x1AEDl0iYfHr4qODKaLS6rS6MKixVfiqzlqbOW8bZMOLpHA09BCzP1JU8ldmNYwhRH0VEIV02fBF
9ox1m7/rW6U69RjOnBUaZ/hUyL9L4U7q73yOzuZmr1WV2Upy73rcOyaNpO46xgCaKbDJAQj7frrB
toudSPwU5qJHsmlpwxYrZk6Kv8kKrtiXAAI5vdIpOzdBvVwGW7Roc04pKlK019OK/sdeK9V2/gUw
4xbh6zTSFfihBHD1peT9fGbRjmRC0DLBqEfRkU9qsGp4TgvlnBXgUjfv3AGlHEdHDWaLr1Zhw7cv
LAkmUZ3mAgyw3jyeFxN+JseKO5rzozqAJng7Kz0zYlJNMnOCMwLX49pnOztIgFwWEnhLs/Z7USd2
ztboypgNQ1RAjVqMqQUksOvSW6981dhIIkqv+1Ex8YvwJt8eYaOUUF9+8FyQdvUVpE5Lr4oEuhM2
UcSUoP5M6Xbta6EAcS2mBMgeaAjjtBkl6mpCMB892tV5HK++3BkRWje2c+e9XPKxX8+SXzXZq/o1
t5cIbeZPaeXQ/nCQ4K3PR8Vcd/u/fIP84Jxyjr7GQlBJI3Bng3cHw7wATJ8r4SBHMAtMuLHWNsKB
RKeC1vTou/Jas3RoUib9U4iZCmvaGzk20JHMDJNQM/X3kRCrngNNf6pOv8Rz3zDM5XPsFR1xlQ7Q
k2p28C4MVq+QJ68F/672ePFZJwy3MNB95/wu2eKyYGG6uqGf1KFh9XbyFIbniKRF066Mf5WzzXnP
hjv+uT1oN7WXrUCUqo60wGbKtJKF0xh8t+MNTQfMJHI1WqZyEAOdQvlUImRcu0ClqjI1E4RHU/Pl
nQVCWj2p9vU93BJCY0spUThlTW6X3+5isyF4cXyWZsWXkV++qdzFghaMbOcS8I+YFGYfTxsAQZym
j17eB/EuybULJqZ8FpDhwPx0GNGy1jBmoN7jhAhVcF/A4TQ2ydlMiVRvrX+HrMKXEDhuZyjZSgyr
8LKFKjTiXIrA/bS9xc64Q3xaTRKRII+cSo0Ub5eqeHom+X0qrxhdBA2NQFhyl5ip9hcie+0Nh7E0
bVEz/J3+jmgS76peobewagkkgNKjMVRVxHfGZQFmGPDZk5a0ovjybx5eGpD2Jp84rAoNnaIRD8Wh
nV1hjpq6pMhyfQGuVTrXwgJkf2C3DCHCs15K9qtEqYjXDb+0yJDB6jj+6KPaf/xOzCvSHpyN8hsf
S8z8h9DN3pQme9YRehbY6hiNvyc6f9MqXTTlRqeXxzLELYZUVqJQlLG+1yb45xSDyDPKbPHa9AfI
sn8Txx7zVnoqs7F/AHbgAXTVDi9kaAIIwWDSBeOMDGxwpfT3XMFqXdR6b/Bokofq7EdWTySsEyih
N2i4YAakxruNLHtPz9aVm8eGmO3qumKv1nXmtnqTWbGCCSUquyzfuw2XugB+AghpHZjchf0rwP2L
S/go99yoVy+QZ5EaBlKHP6eF4cyk1Xwmt9BLiExcCLWfJ70Vep7pCc5iBKTmTS3SBtfr9AbD5JEk
GbYVQg+SCuXukcvrEoPxguE2If/BPJ8OCmcAi072fLQS+4/h2Bgb/H2plNYVRvap8XvXgIXHMTqR
gyZbj+GsqcJ47FpLlT6uG/Jf6keVPvbFTse+Pt7vjpuAoCe/h7r7h24tUgCCnQkgkVLTqAUIy2Nd
NrUOHyt3spjVNVJ+574aoaa/opMqKFJguatKHRN2cfk0vHi5iPJuauOaRzY7kwQlXzPzwJYBzkSE
H6+SmXFnFvYL1vUSFsyrvECCL2rKMcn6Tcer7YZqJ3xUDNdMap37Czhy5yg/SLMTdzUd1FgGM+4I
Fdr2ox5Qv8NWOFxDg/0Jt34FZ+acBZHFg6NvQxz3+oR+CPlQMu3ZB51z3eO4vHOCQygPKxqVF73m
Uz2eXpb6ikWloYiZZElc38qGtPwBiGx6BeCzmdJyejiEEEETWav0KfF/r0w0ylH1kDME5G2wkWhP
3pD0Ed5NIg4Q6/FIL6nKfSHAp/tiAGnNMd1/3C/NrPJMJ/u1KgZeg7eLO4fvfmj5l/q3MZF6LboX
EPcrYtrun/vsduzg0cPJeNWpLu2w0e6XQBbH/0Be4pv5bMaiGa7HTSbwPKRn58422pzlzhiFpWtp
3PqIdwzPAINNFHD5VobDgpWr4rTtcQH+WMRJC5HpNf75gk8rwD86hoXfTXf4Sy2ksizM8J14CJmD
4IXZpePq5w9xEEH1ZUsIwvWn3IRiNONxa8hlfrHGqMaCjinrlamQKamWDTYEu8fw54n39KTpT9uy
P32xEZ/3lX4O136yGpK71wFzOnmtBVQPJ1N66aZXuhkXcp6jGTQDC9o7IlZOg+Y8p4ZFnbZrWzBM
2eX5ef0IzUhp5rvN0cwE4QxzdNVVOaOJN+WLMARonBGOPlIAgS1CX5MbXBwhQW08EQ7xwVZ/ECTv
YwG2SoVT7MZvaPtgkWeOdmEC18hAhOyYZ6uH/Dw1qVaUBfaWgdgQdN1AFLoen81D9JzVYvtThLr6
wtyKYtM4z+yauRsmEBO4XVE8lUNARPAxqrdgHHz3Y4a57PP7PmCm0VF72P5/3/TqpneEs0GZpXyt
W+d2XfA/Xsbs/fiivFzgcupDAZv+biCNr5752CsyjfTsVz0R07zPMsz6llZJi+Wp/GnJP4bmowte
J1bs3s+YnKhOjFC1cLxVgndMZ2JgDca+PICBTVrEOhWZVDIFOAch+jlcWWzdKHvYVCCijemW92vr
iuIa6Awf52gmX1hjhth7K9r129eKdHveU4/o5AodvQxf8o6e7Z6+4JbFIK9wubdygNllIHzL9KeN
uJY8mAbzyT0bOQjCBDo6l8e29C1SXhySqE3Ku81j+xXFEIqe5AgcMJHE39hTUbHqwasKzLd/5C+z
5c7rCinFBaNWXGFqtcxDsq038M6e0f2dH7ROL4YzK3jgxgFK5Gh52Q4lc6lGoOQd/Nx17AGhIOTu
+NJ4+XLZWVM1bVEg88tN2UZUeaJTp9x52AKFLL5yINL5hZ1r55M2oPaOTF1P1TXIrwzumAWaHqgj
n00b4NVR1VnbKy9lUedIutD1hJ7vCMeojx/9xnFxhX5wxOmhSu8efkZf6v9tfFecILNmKwy7MgKz
eeM5g7UHAe8ISnVRLthUtcVhp0BE9Ca18moqtE5pq5qcbBQAbKSgOelZ3Q2HrZEInIbuWaChYRiy
j5iJj/aYN6fbbxpxxEaZ0EnyTt9klc6xi2TaaV9Q47qV5TsOS2zlFj8862VybgXgu1J8cki20oKr
H2w2fdtzhCFGN12l9KtfSE6IZPNwbYoCaVzI0qp0vfEYUvXiMlAQDe9POrY7eCnFWGQ1c33cYkbv
sKzQfwGD5E4p40vvb2b3dkDpaQYDWeE/nomin9pmLuyJ9AWZmwjNVKZTLzLxK8QTH3ofO9ams2Ru
xd4KbxyvxrhYddx+MbzQKdL7Xq26KxLPr+GRIoo5j0Alw5dcemJh0q1MZTXklDUkDthfZBt+r1+Z
2zIgi9e1DsC2OccJr8HwFYAj439fefFoKdJfG4Wv8ROitYthwwgLyMoVnYZcMEZCjJAz+R/59WBY
RwHoSrI0my6AY/oTPH0FvBq7hMmVDB3dGRqqnesX0/LsZEWBVOHR1g2SlhtUMKz1XxSV1dxcSqUT
1tlJ5yrtHIU8dtycA50CA+9I4Q0K/DzuRitsyhhw0IBYElBLDx0Zp/8PFiWxj1H3eNMGLzlVlVX4
V65qUPksYVuybahqHLKBZLMUALZ04jXuXap+tABuUiCG7hFoMZe8p5ELsvXXhFjuStgFbsPgAZvt
58vnFt/ZBFnnLAkGcINAVoZP3bjHgjKkIC4K9HDGC3YyFXhCAnLJ9zONnRZjLRF4dRMrtN+sWJMe
6gUNv6KGDiV6DG8JEaP47B4KZMqQTE2CxzyeVN40qUj6FJabu4kLJ7CZi1M4nV1KyhkGuvIdo5Lg
ThFEsSQeYfkdiWBvilKC1DTDgvbO4EAEfEcibeICleIDq2zXGSB7h13B8/NkwLxl1AWZVfSeh6vM
s1Om+pxi1CLBncfqGAKN2rYKGjId7FKMpT7RNKIbKs+GCus5Jrup/1pb7h63OWk/hPdu4OW7l3f9
8G//bByl1E7OEsjULQmzSfYPTjO+cOJcRUXJqJbBg6CK4Lsualx4ZXVCnVayUas9yiiTbjT0StCc
TLNOirYbohmL4fJGjRGt6lRnfbymZ/gaFuWFlgdxFhb409WSiTBSIOlbDw1Okc5WPProlqZuJJVj
fu9D8lRrnFBw8FXF1T0PaMvd1UxHmAow7YNGFwAUo/iyg0KklszR0/yL20OJyCBv7KImIqevBCwx
g8d3MyHqy7f5lv6UhgF23mDtK6nZXUU/TULFpEE2hhhLDr9ZKTaDnJHM86Rvs4A9O0ieCoz/uXjU
BKd9j3rHZtKzwCHzIp1NZTFFLjAuD/L4nGfnBBQzGcPgqlFmXH6Gjta4G0J2z+ehrAr2cKP9SHqq
Es0Omm2UsHDNC3ZU0to7Jjp+gxuzdjDen8VtU/8enMSVsoU4+DcKFgOEgYmPChUb/SLfS1NpSNjQ
ln6rvCmfzDTcTGI5I78/QwNWxvcISCe4hg17e0HHBCUJ2o+iBg4xDYDUymVn19fRx1oNK4oWQ0R5
HgNm/IGtehzfTyZEi9Xe2DDvKglHbygeAH6XwVVqmohMmLUpaVDn27teLy4DCSjtYeHvCTqem5np
qCY9wqPRqxU86bVmYEkh4qnGw/lRayeRXGB/kJjlUXuNQ4oPpROGsyKVxlHZb3DmxrdXvLBsmA8y
7ycPhacNcP5v1ve0VwGcSDp5Z8dYTHiDcCY+OoYoE95yYnNNTaF/5cD1C6PP5yobaC9oD68QLCAD
lu2ylzqCxPqK3kCSDop7hGgw8fauvTNwE/pEYxauA522/+TftgoKjmbFZb3td4Q4mHC8uoU8Kyis
fPdyS0rLOiPcf2/1dNInAo7DYso91nnsaMhLyoVOWiz4mf2TwvRa5gPBHABy+lzM0RPquYuDxQyC
sy9LTeAq6ZddWFLLcTD+rQsv4oldkRnyYabm0V4qtmREdR6DGkISvxqCDPe9ryHb9D2W9WwPdih0
as6BoF7UjQ6c9/GNmHTuf8FUEekIwMYZoSdU3MnF0GXBVLTL9IBBcC6j28czMrQTCCHLDfZWm4Dr
vAj98nCSXEpV3wasfBWVb8jdoLBmRHPbAWigSzekVBpChcCOn53rS8vhaACe0LVwv7UmfWeGyDLI
BbvuU/TEyo16HgLflYHb9Wfb7eLxa8sLNKW+G2rA+dHXWeCjKE9k+3rGnthEb477YVGmXbINQTqc
S/ZBUZMII+yqEUpCDBUxc3xCDpFrIUWzC7awIkdvC3AayEbvDwevceqkmwPe7ID4Hngv44YpLObn
N2YaevsdynExSgAKyxUnutUzRWMnb4gU1O6OUW9CbBFN4xoja9voL66CINXRwFL9lKTepWCXgjoJ
U1kqHkxjQW2WeMEFRbNFaM1y56pR2b0R4LZX1RGZ0PRD7vweNLwIqstAkJDNlUQu6PPE0i7s1wv7
327oNaXy/pOxGlBW9ohEy2/yEx3wCGqDp+NsUr/nFik8yA+sloCDwjVaXLzfH784olqfiFtwi0WK
n7H5wEvu/HpEQHgVQ/Xo2H/WWiFXcjw7KuSTSyG/y8OaSfuJMvLZIr5D6wedGzJ7PKCYLcuU1bh3
pi3thTEJ/e7shB0CtC0ulwH8Sg2DHxAFRZxArSJBhRFcDOBLGfGsPWZu9I4nkG8OLnOxdmL0bkob
zV66Qjn1TR3ebhUZmuQN5WmaVfePAOyhs3hYZaPCNNmbNn2Y0HuaT50ZaYnyvTNKreQYxcfhIG+F
DxtaAbpOWYPqQFVuSGTVxQaxA3b4MC9uvsPZoQRvNlKkhsWpo/4o2Uyyi5pSKAO+plxiFv/nWL7h
Vl/q4Wv/NBpdxC6t1UwV5N8DDTqsoXFoLQOYc/V3P928+XGynRHnf3TksxZPqlVtnbKuVuqT8jyf
zUvzjUbsk6VWolnEMSLWuDbkYl/nrf2vopo0WzYdckIF2frniUsooXpFd/7pafJ5Wry+gBU1T8nm
CJ6GHUqeZyQkfzbZQF22GxFz9/SFrLMwrjMhHIK4M3IQQtu1Y0hVso3B6QYtWEfHJpwYbxoI0vmr
ojxGK4X6e9PMoe/v7Z7qen/c7b5a8nDItF1iAVwuP0dFyTDmXkC638S11p6VmCkG3qAiZbDFGswu
55bhmYUR9hYNKNlxVG0c7MjCCT41bICP0aaAyVO1ouwxK5cDH2pRyyyYcsZJLZfFKrrbvQHUkpOC
JitSP/UWjaN/LTNQxZZOsS0ZydOVAUatQkGzPNIbrHg9ISGbWuwzlVRj97GNdQMSCuZvV+hvu+HX
uAiJzVUxbAaN97NChkZqQkoSygKsgfhAoWOKHyOnH/BWM/S2nOhaL1QmQp2/U/mfkNx0YSoSe0zL
mW4a+YzgRiqt9YOt9jGZf551+GYtYwtWGzupi0zjprF8IB+F2dEvbW0M4R5RoCVnG65nzPJTXPTG
2LZIu2dUqPZNRe6dhX+OtHXXlPlf8fS5sy6bcvb6isHR73K8DL5wLIe5T9PWPy4otPBQNLzChIgO
9Anm4AjTY/3dQitCpSTSGh478R7Yy2VB9zJpVHk74oVggQuMVA7KpzDh/gXko+SJX6DUGclqVhyS
YvRppIJtfVFuAFWkNmfNwrBBrSGwYalErwM8vtmqJxQ7ik+hDSn8zH+58Ft3TH3wvwKSpOcthiKY
CCk+cGgTxA3jLIq6IeL5Wkch5+xnt3zBwRL4YlfTHmH33HpT11j5VXctpfscsDkv1XpzJeQ1AZ2c
qY1vuGGmW3pfstAmqwTXmwa/BH6KyvXZSeLfihpCkAgdK1H4iJSU9ftP8hStIOfAlaBnjVOQSkZo
N+KmT8s8vU1LQJaMHad3Jr11xd+/V5PqVDwwZzBlhHng2V2JaSE018xxNBsNm1Wq5evd259JP7FQ
wHRc2uif9Qb5mCvK33Cq2BaIvgvOGHvaMYo9TR7MrDV1ayXZijeQTvSrGXRn9gu8tB7iV73PzWha
MCVJl77nkcfQVX3ZcxUnAvqxyuXUdCKVozEOpjFWmV/Aq8KmH0fZtPUusxneUzdnFTQBgkuuMEp0
/N7ieDT+/NE3nDjb5GO1nrPJCTNPo1oSDsZNkWNfiSSVe6nXGqGMGVUjRXtOFtIVxdOmoQk+VStZ
2UBSofgMvo/1u2pH2b4QIAVpNTJtpPWdHGMU4Nb+1swxPUIjrNp95RErv9jCi1uKoBUjNHbxxhDC
s5Mw7p8GRbJwTOcU4ZrbUQfY0wiOQWk7ZvAtIaZkWqmSjgDUDFBdjcqlWmttnH1NTdwNl+h6lO/c
3ZQUWps2rYLaEWcGS4PFf7f7T8JJYF377Md8UBvAxtOv2ZPpqVeBcNnM5VdfcutGPDcwdd3QqIJ/
WGfR0Xu5slqasvrbqHQKF1mYk9JyNqY8VZ+//llTY6A3ESl3qe+56ZPsWm2B4rGJovmw+PGiEWFf
DAtEKfYxoeYFif+9amq/RRBtQPZbiYTsTgFUQIOSKWsYe3tBwjPlqVdDv+j3Rg12st4WGw8uwMLr
L4ynh/5EODrwzASJkcebiNtPEHwwRnj7lLz9WcdwmCIzEuaNylVAxOQQ2fmlCU9KKcVq0g2dssJv
YJHCCVOx0Nbi0EYG9mPx3JeAcLetTmQbJKzSGfxEEXNM52Ai/HJvsBIcnVE93XO3O/91aLp7YcvZ
nEGFXiMlFVWP9YxacTfbto89eHhocjq+fEtl9D86jZO0JkpLFo9+gRA7ZvRqNm61pIbFKh5HIhKD
0ZNtFPki9PaliLuw7o4n//3sKGNDeQVgFc6DBuDXavM1OKG2FzB4iOMs2Sazc3ad1qiqmF9SXzTu
evsMASiPGm62K8DO+1itFqcC05ZnX2cUZtvxl3rvEowCwI3+YciiN0AD1tCu0dCqHhp0Rq/N/3Mg
+nzzsfhicbFYm95wGT0EJ8cYyEgRh7YPb/p8WiMZWyKb6GPv/4zS/hWvAbM7YYOWGmVDfSBLNTjs
Fb54bQWqGh/g/PUbbgbBQzI9IXRvqawUWXUnPcw/z9YHldGKvzL2DhNRNFzpnNbtOF/+XcHViQPA
AiMbMynEsY2+kmcNQDkBQWCE7Dk0F8JlGk7U0giI69wYbmlVx6TNjgUknKzmRpN43+ihOmMt8Fiz
sh0f+BiDZldk9g5o3dEjes7tX77sMf0W3HaDCdh+s9Wo3/P/orzU8cmU/XCTEIGS9IKxuwCJftaw
TcMF30Z80eJQtPevBxyVGuks1XLAi2AQYaKUN4mPitwL7/UpjfqpNd+YBDdPYOtqjl+qUtGcl5y+
2rW6A8UiKAZ4DsUUzaO7Gg4U3IHcD2MV+eJaZmw4+90B9Crfle1jY8GZu1WziWVxwh5sLzmtswgN
TgLmghC9J8zjT2i3FEsP8kSfjmDwu4SnHKgpMKWqO8BsfyK86vcN17gHvbMv7vOmgJh0vnYhP5RI
FVN6IVXLiF9QGvcsd61NaxC7yj09cGR+HYogYGH9H7z1dA4TSskIHZGUXKmnQr/Ysa7NpZIcm9KZ
tt2A9FW9EyZHXdO4a21qLdon0bUchP0WpJhqvGpxMS/IJZDqSF2bx7A10vjqgOQdOiXxgsFA/Dzl
7QuRm/DOf4prIpZtB+nHCIao0EBNlX0NkUPecHJ7zhJbT6KX11Nvv+w4bxOaWhxoS+ol05iADWP5
tJc94pd1YCsI+RadXXqX3Iosvpi9kotVnqjppJn+JXGtSqYhAsE3eZQONcmTwiC5/7JZ6aiw9u0n
jh51V5JPiZu0Kb620yZVbCBsvEsmo3FqiiIkAB1U/jTwkyzXkeSWhqpE8ayZs6VTliwMejGLIp7o
nsB5SxsJQkAbeTwaOMJS03WwsyUWQWYjiy5ER22OBx13PP+Sjx+HCMuscRAF1kmrgJMImyHhRkH7
x6WFoTZ4GuSeRg6aSkFmxNT1qQe4+FVaYGGCrF8vD0/eZCTC303wkL4FCYB9hHHmhYtamaj7B5sv
NIwPsQFBQWH9JfXbr5h5Fzm4dHfiHPgR+AELy52kM27M2972KHTtxhKEFzMDrwxQY+lULZHPKYdb
2ZrLM+UAdGZN84o+LE40j2gsn5KMYiTPcgEAsLZy2J69ySiNv3yz+La5JA8dfCoQ5ZahWJ/5Ey0E
7Ggn7+2hWkhWCXb5nBWFy7/Ql9b9ey9UtmOi0S8BmaNTYn8/WUa/FijOKSnsJx7t8qPGBnnNCQDp
YXRrQEafuf8mSyaikYHhSx1T6pNRPBvdcKOr3MSKCrfkbs9XLUCOgSH0+3IQVX6C//eg7aZMP3DF
KqIIZ69wItmz93kMrnidDeXDxDIr0zCPg1yh0IIsE2+CwzNpCwZdUEKHWBK0TkaHbHOHB9arQcWe
rZ+PHM7DTf/n8z7cLb2NESLpJ+8wfOEFntsQvZB0z7U/kPsR+LET3GnYgvs01ck4kYa2pTjBAMjW
0s3oDb18tT83V0g4JOr+gPgZ1GkMS9RK87hQLXhbvvdZmXRdIa6mh8aBvy7QWjUKWx2MsEBeqYOb
kabzO2/Uh/6hLqUr12Z0wbcb+PyhZOfXIT8XU5nBjfwZ93nve12TeMhfTSMKHZfFHrOjaO7vSc0E
wTJh541k4juCz2NZLXdYXfT5nhs/oakV6GvVXqEcNezDXLu8BR1XCsMRX5LTWsdU58elmyzh1SOL
4dZ3n+CCaR3Ank3Z0QqmHXuiph3VYUCi2PGggQMIl2qrcOtbNoSdqPq7lsZNoEgOGsufiH/ob4Ge
TxwEOPy8EyM5F8LQAoAAT83eVTvgUCBVizXVDPxJQSgsHVVwe28EboTqwws/WXimFjGMC6RCtffx
3aBqdx3wQiQqtrhJDUxIBuFI2c9oGkxnIWfShKugBpv45laTi4gxHzZXgBUjiuLZ3rx016AnrmRs
JF7BZZWOeqIKS/lXce3RLU0mGLUICbCMuGdh0lxIcu4G6yzG8+7gnRjxQytbVWtSFD+5B2d6C+ja
A+DTQEYNdCnLVkt5luMt0/YrsY+jCyYcn/Mdwp4ubLH0gJZG0a2+nLElQXtyHHcnUcU3TndwUJG0
nLqivLBeT22N0KjvP0mkGYBi0mJ4qpf3fXmDwc6oJyawXv7WP1ebsQTi36PoseMDlAYUgYrJGWuu
WZ4DzQMRqbQwN0wGU5DKIxbPSwDpEljmq2ZdDo3K4PWkNRc/Z1qwATvJyWDV7JjMyOVvRsg1htif
OWGuk6ddURALSh6GuxazncyuYTqSdlhWC9SRykIFFLpwNiGVy1/0DhXJ8wAC3YjG0mCgvmZpMpe7
1OcP/LDeggThh2QE9OWynaZzHgPJbsJLOw6oQ/YlJBZinS+VV5RhtouskbpJYVm33WnDy84iX/0q
GGgb4PagKLl6LbZNH5tNlzRyM7swiR2XMcrIRI9nMjlSKUPkYMyqq2Hcxhs5JwE++pN/5TTfkTt5
NTM+2hrq5Sqjaenblg1OsEkFqJrJqN5W8FEMKw6FrDgTIABtvylnApvG0C7mmuAHKj74NPV0aIz5
4LMMtFtdLsxK0vfGjMxptTYSS4vv0v4oG7RHJ6I+cJAw50Kr5ExsWZ1VXypqu5SgCmlxujO3A3s5
GuEwMsJGCr6Q25U0qwV1tjg+PPVRwzQPv+AgAzf+5QE6QUqVS/GY9YmLE0FtQXQ3bqLCxTVP2iAl
0KmUo5IXKi2wMirz39Vq/0EmOw/XavN5MSt/xygwPplR2+6aUQakq7nRASdb4wLWrPMH4JeV5y4z
sPySPOaTg7BQQCYAH/GqpsIbKLv78YrbFvI81XWZ3Is/BbUOukYMNdzy+QXcTZzq+YofKgVfsBSa
A6pIx0D2ALoujvheutDexQ1fyb5870xvdF1xEPv3kHcxZr6YELtIA1EA8d6gA2byyJ54lXWwUwJs
voSdTUJEsfHETfqMcLiaAz4QlhnFQ85ZQ5d/rQMWGKG+r2P9IHblxuyXQM9T0j8asl0kxzWmPJEm
wKAYpm0F3zs/bs+bXEEpDKOa4oF13lp02iVqwJmmWr6e04BFlplyAHBgibnSBRTT5iE510yYxi0E
mg+CT6q6LjhIYV54u5JjIHA6stkMACcX0FjaIjrY3jnfV3AVUJHyY5/QLbuMiG6wG0qnU5wT21fZ
BBVnkZuwM6/mHtNnCd/O7nceyLTslga/oh2VdnYukuC5GSWDlcY/ko8be31egqagxC+QJQAtV/sj
uhBWWpmVaNTaJN+RjAMEqif96yXMTtngxY5KgEWLeFOz4kpebCGFcABAliBQ4i0vyC975zBr3kev
/Cy1CzzjFQeHVC1I36fh46e8FGFOlcAQNjgRGLa/vLnD8lJLFyfwldJrUCHxSpWPRu+9Doa9/xCi
AwyXBO0IBMSWnMC7IAuaMiqT6sm8Z9mdc1XnSdso6E522guHWyODn86Ur0GFkMxNHVhF9E5zAp6/
eFxnRW9Xqpc10nlt/RLDzEG0ZtRqBhrTPkAPqvQksaXeq8k+kht/Ut81l6S3It7MGR2OhqL8Fkgd
M/wJThJolBMgGJvnDp5A0q9aqxTJxr4tB5r0F2XjJ+TqsXTLFY4FlNS+xA8jx6mDdP8PFdD8IIZs
lbd8SGRLGUMs7asTdX9UJzVV7kzyKcr7m8XlqoHTNLk7YEaJ984vglGNm7EP6s1cGjBkZ7ZY3y0f
MhY4aX30Lf+scRGEywPjN6VjSAJfbcbVeaeXOHUkEk15BHpZSff05g4EShc9FnwNKYWmb/mIp2OI
h3mSz1fqXTE3xhwODjFpiC4dG+xUSWapHAHubpwMY02dzUpo6GymJt4RAGpYMgpA0Cp/ZouloA8X
6W4rnyJM9Q5rlJe2rEkCkd99fb+Qa2yps9k8c71vMJS+QVS7wO9FO3PuhgQnU20NgC3F7PeXG0nm
g2d/eg==
`pragma protect end_protected
