// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:26:04 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
o0jFWHhgpJ9GDj/U638PPFNoRKzk/9TOGzL3N1MawtNRhQsDBaC219jWBvxWviTO
JO8T+Z3zOGp3GG+67XLF5L9xdKPUeuHADNf4brdJ2DJYhpQelKKFXf6kPPSiwozU
r7f5uU8uO4yq1vBBFqq7Rij6wb+43Iu1+1B8OSPhVtM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24912)
txqcQLAYIwai8n3XGgNF3MTcnIPCvffgKQdkc/7hmu/Ky75pYPBwN0ufStHaW672
G8r9zzgCt5q/joDAbKFFFgYK0TUMi/MXqHR6XwJKZp5ifm2oqNnwM3ujTMtOuOio
AXJwc5LsdoeAxB2Jt+B3TBdbc13Mp0D7YsiWLiKle788jXH0fZy27aV9dzDsc1bB
y5r61TgX0tImn+9GjlIIh3u5S5+kPfiynreHHyJWfWB+IpjJ4PMtLjdFuGtXx512
m4d40YNjQ0u2VVWgYdoxuxPgn6aJXPl+nmYd8tuJcaymmozTE+s7wmakTfcgz09/
mQI398qLOwaax7lvOLo/2e6swXvEafYHMoj92M5WTCKfFw1HfK8g5AdVWq2bFem4
KFJP5vIC6OdsyHTiuzeK1lC5eTeDy+oSEOfmJRCcppUj8F7yG3JYGJ+AqVMvitfP
4ri8guIpy+joM84Lrfoe1cjj7TuhTCOeMAwS+dsWQGsoeuA59RUluOjUKVid95N9
A+j+h4Zx0satx9FVa0FfssTkEReu8c2ta7ezduZazu3oqGm50+gtihbXmtprPks0
C+pxc+wANRWzXtQFWrOYZPEWSBmuUBcwL6SZHhq7quBE7KWvfQ5se0pXQ+OwrVsF
39Hhg30wLQOJO8ugaz1uRrmSZc5vAZBvU3IHfVQ/mygL+L/BbYF5TdfqV35Mbh8V
qmaiYGSbiQMA/NHPEKO3684Km6IJGytX1stb42bBtVaIhIcg0EbXq326PfIzP8WI
4X+LUmNPFo0LpvZ3MpPgSGFnewN2BSjaEm2p90i5hsjeTfxj5/Omak8VJj5H55jE
11qt4tIBVmmslag2bvVHeGEnPfC46KaevmT/zJnrCr8fjBrNjEZvMmmuKNy7kiaO
bslaSMJXdJ3uP4korfSH0CN5/G+nEZ20kymv60DO0PRgWQTz2pr9RjhscOS57NaJ
JXieh25Wy2JA4UenDhshApU26i7bK/1jYtEbJUJvVpB611hdNlA6sPXcTyhU+p6y
jTBuB0qpXPn5ZAG9uZc5NoDzNRfF+rueSrLKWGmPXrdfT8a+iwt+Vlzbp1Hf3j1E
pcsRWwfynqEq3KfVYTIA1iULBF8R22DE2iyzbIA80qerncLDp4do1RdMt/sXzqUF
2wk9SBJRnCWb+KORs5u3CtHH3H4kUpXXrRJBshqZcEQ2NkrpN5klZK3eIkx0x75w
pwNQnMvdNLi6URK2XT0KHEQhdRWx5TIVLEn5Ll7Kdz4B7XdvO41ZeY10Sxavubq1
IZaWARu7XnXQ7cEaTG2m/6FFJWkJ+wMZKo19GUNZ7gqaUxf9iljkLWMnlwUi3vvS
g9Akn0Tmz4eax5SqiTZ8WLUpBOBL4OcYliFOyiZTb7aTMOFOyiZ9Zu+er60/C/Ke
mqsTomV+h6ZM5bazoMZOIp/7ajhCBZ2pNp1Sbsanc+6IABVeKPQMw4S6td02c54w
ZPS7eG/4sWEkww30h9gv9VeBGZtB/RweOZgtxpxtXWNGGfr0hNKfvCQ2VNiYrCqT
/NMCCRss46buaH7wOPly9Hmv1yWE2jVsjHqdVYpEolW8vg44bx4MrERBrYzmeVOM
gRR6QpoF8twnbky2hasJdzNCXssdOFtUs7+bFZdXz6vVGRcNLeqWjQmoNZljkoBe
bYMXgP2dugxgbSg7PzytU5e7VEtxvTCkfOtmzg8+Bw2lUyteg6sf89ZlKJTyKFIJ
akf0RLuovuFZ6iCgmTKj1Ro8HYo111UxzciYtxJouF0cVq7qiIPf4JL0XwSkLMq2
RrmtvcQP2y2/mwOkZSw7WJa15O2ZVlhfmf1+B/A7wWOMZNTuHuYSpJrMV+77+kNi
GefceBVY4gX34gnN+NaavON+e2CUVRYeeOZ8EPX5gjNk3YDO2g6LqMQNGd0cdQG+
8lHRnfbvXfLVuaoEoVTlMdwcnv7hT+ke2IQ6iwg8C3kR4LvuNprusmwvWEtPkz6U
siEB9zbtzSB7D6gNqMJ2P7POV2ZNEMuaTt0Lr6x3tQYyPmb1L7GkHiboAuoAbmnB
jmCG1Lhv5TR5vd1Ab+TIVf8O1rcQritPGcUaUEPn5kS5aJW8ZFq8mXmMl76bdoe1
NAjoPwvW/6EXTTDKYYdYPNHSvSSTKq1qG+2yhs3EPsPf+x6+qKfDTMaI/Hd7kpVW
Uy2sGoTd71BL7APosaHONpyqwf9LwwNGcRNtg5UNNqd2pCUSab6DwTybaiWRkzKc
AXnyUfrwm2IyHDD6E3FoE/xlRhHj5q2S9gWXfWQ+fqm6moR/UwisN9sOcUfdIFdt
EujBDMXCRYwqM1/1T5Vr4RefYt9t3lD12fhGPecqQXPTId+2v2ly0WLh9o6wkeSE
KbUgvrPevhPgbW31YhxTp2zRF7g/Tisg150eL6tGMhQmnAUerI/l3Fj7sGIh1RCp
hMcfb1xUEEFpFEkcqyLDTmrBtNVKUrkXr09zEujrK0x2Q2T7O0tMn6hhT6OPU5Sc
K1oHd4xC78dqiHRbIUyHFLHx87oA7jfrt2Hzenvf0XXs84cpvjrm8vokbRJHOYYt
ANGCWaGnhY92ya5/9X+0WpJUldp//F89oDGq8zjsxf4xma4jgTcjbFBEtqjePtRT
5Ul50hvLZvvHn6IuUfcUwUJQZoL+xm4L4pZ3mirMmMDgrtw+ED9NK6i7t4bBYxJQ
wFDxOsuI2/CHHnv4tBaUvPjSD5REZea+I8aowQwcJ+fJ6Zc1vKA6HT/DBwEfZXd4
SsycAk9VGeDPdSmDLPePRZT4eRQS2gdMTJE+4ZvLyAkIxaCXCFDrDJyq/lYewbaN
SUwBtPqx3jud9UcT0Jd4nE8zT40UX9JPS1V5FIkQB6vs/JixMWhfXxw+IYQLQc0a
A90Mi/X9feHuQgpXJt0rXU5vgjl+whYCXnUokcn66SJeO86aSRPyCnV8SRocqJl1
033rbPzRQmv3+GBOxkSUa/SSulNaOIDmj1VPMbBY3Z1sOmrMk36fvXb+q5+fLbKl
tBQkQmHlihP9jTo4i/7gV3rUG9UZKUPh8E0FfGztmfraTLHOeF4qXm2PKA47JF86
c+N9GPCNia5TqKFl9GVs2RHB+nQ0RlAzaeG73slNuXtELOFSsAoErfvqw3YIvLLW
fvXAdrDHF2WGmDMxJvyGizOGz7pFzDUxDEyxAZ8k4YBB2H+uE3NzftalxbVQMj6m
E95fpXf9yVHv6mPwJzYna+jMhwxefAxx4sRKAP12iKwG5JprG0OJgA/g47YRUzTP
D3N22uRlytqF0XKUZ09k18QZqhcTs1iPgncLHi9cQOcxSXc3hPOhLN9wIVoqx8Jm
v6G6yJhxnosvoPvivqowcFZ02Fbf0u2vtRBStImAPHrq6BxSkxziFRpLPGpX2Bn7
bNide/YFlu24mYojoaXvQpOQqNFL0uC8Os1iyMCVQqbteLmKyrGACd11x4RhG50R
ad+KIcPdWsDtiE3+ncsRZUJlgiCI7lbX/ifMCP80Jd1+5CG+dMrYLUIrcJR08AZL
Bwc/DnIEnzCA5DwVa7I8+HtpLEHG/KwiVGto6yTmssBMZW7KXa3oQH1NDhUrVOHi
w2qDdAZoxzdtNcmIkLkwrIVQaAbihMhVOFr16LB8d1EslfKodQgJLOF6z3IXZdAB
/MiVxB0iMiJn7kmHRiDz+JnxiG5m3bHn+JkVHpbRJCvg6EaKHo1ZZ1200WlOx/yO
36hnabvivBq5xcvD7qkvJwSVqLr+0t+BZGV7KUfllp8XgdFrZm/FMeuFH8ik49R2
BcDmgm3lOWzYUpSyzhepIVA6SHt17dD2TdGsG+nDcPsORWiOxDF65ZZmit6T/j0h
hjMpChaKElupP/3wlT3ckJgRg9RhjjkOlVct4IhRe6DnSkWUvBksRagBEBkhjTcN
xF9KjYAP8FYzgrHC//Od79L7kyDvBDwfieu8twyL5DbbtygYjJWOFnIlhR1qWVkT
1nkiMOh+T7dY2dl3QWOEwrGkQJobtr9NS3KBpt3ttz9D5IU8owAPo9Tgiqg4tUYj
1tU4xvP6Gdcz1RdLhueV4iuy5jK5hOJFO4OIcXQTOv2kIkr+VhIIR6tyxgsTKjmV
LyihGSJZlR4gR5wQLYwKYJRfsh9v24lNf5QVl0vuWl6T7rIFVGDf7fsHv2biAyXH
qWq1+9cSPqUom/FU4dderQtfX8AAHX1tzf7gmgYQV2nxQ2I67CqsiSJcFeMIadNJ
vVDOsnP2Kk4zPRQnY849xW0kEva6w8pxkkY0478lAXp2bx/hwZbs0QbqBVpg0flB
bDJsF5l8vv+YiC58+ySUZrBoqztRHeUsolJNh7BFuk9kquylwUHXz13JSSyIYWgP
PkUfIA0gGWhH2ayFjld7Qua0J/H7B3gn74W8VUrH2nwX7WLPhi1jLyb7bDDZVX0m
dYR/fvRLTISdeeOWav2YFeaMSDrtUlxQDfXjj2M2Th8n4NX+yczfZ8E5Qh+4LodO
sHy5VVN0srnIQQH5KtNV+qoF0Zmj+qWxwJzzHQQoAX0fTH9kZnJ64fWAFi72vb7j
RGqwqDfdiG+s6Ijgng2wL2ICA1xT78yxBs1tEl+Ua7DzjXxX7Ba2YhFJQSGqaqXQ
mLiUKU8mLdwx5GN0BnS83MeW1ckc8PvHxZ2fUKFuCjWkyxqyD8umhlvAnbwgFlVo
kjDk1Jzs7hoAehvUiWRl/cnnuG8Vz3D85E6nwlNNbBocFlzjlT0/e2EFOhBUZ+tV
JVJNQdL33FN/NX8oeXDZzSFjkXa4bRebwDYMHvEdND8ADvJErjj8ifAyNt4NO0rD
38SCbSR23nLrWQYE8GiZbXIjFsXeQgOkdWWHGFKoz5VvlVL/g4y3yLcPgzGG2qn3
fh4GspHxYOKbN/OachheE1vHGsMgqkchupBc1Rz/7cFbK5CsoJ3Br2zcL+pK3QBh
YNVjPOGl0gTZKhNnMqH5fVJmDTK6Nd/SxzxmFNpQfgsz8dtUPq5l5bQVmDJV1mJk
HUm5XlkZfw+Y801PQ35oO1tF75TjFXSquusxHmvXrIznRpXeAUzF1GyGR0ZHKat/
7fj32jb6yHJePTITvCIH0tRMFwaT+wf2XNm8vtDTH3MXf0NPQE2Pevz0B5xW7F6N
+IUXvS0KmtlmNZsH8rFGaAQKS+D/xv76VIj9ofxFaCKWXALue2vwLJ6N1B9K+XCy
yNE7v7pWp8kveT/QLtXdBpfEkZrtNsJR9AafZuscybPGtX1B042G81DJy3WzjyyX
vy5DX7qebCPkwFlieqS7KQyTOa/VGMgdyRMgZFTBNvsoN5XXJcHgFZz3kzQcPlKb
58CPG1IYW4am+lXIXObR6PNkdnGvKKM5skq04pBsKYerH/Or3189YU70OhgnF8WY
61zsIQEU/bF/j+91qsHUX3n1fJ4Hpp2KH1pQ9pjF3VpXdqE0vyMzSD6yZOupCrkV
P4jg09M8AEjL6p2GkPAth2QOEf4IHXteJZdFlKtAC9+QReLaAeTGzLiO+cG1YZ0w
CaVvAK3zvPO/ZGT8mzDcxvGcnK0zzLfG+sRHzjtxIurbXfg1KJHpU7FyD/EdIg5p
NW803NxrNPNNCCCxmGYYohfA09+q2s7Ecp3+hIQg3XXxr/KMkP0auTB3wDO2sJf0
GS7Xn42O3SF2KaBCEMVkVpzK30inc4ph21C0jzzKM5J7orB+5QxAc2TlnIIA2by9
9Eo6BTI8mMSBpgL212G5pKKNAX+I0oFqQ50pu1RlK/OtNXl0sI0TLZFLKQcuepML
d15UuMgWIx/QKHamowDpMzlWnhTR1aY07P+RHzPOG5ca3RV5lXahrjNeDDerY50l
288H8vfIbklnyvtMutw/f3u5GwzT/wxgBb6wobKRIKpE73OuxPaMek23B9NZZ5Al
/gj43BcBy8upE/8i8ClmsIHkJH7dsjs87DAcE+lcmkcOFRkmmjds1id22x4BvmQ2
3LA0e5BQ6Rw63tdDjke/9FwgMqJc/0gOw04PjU0qf+Rj6G4jL1WpdXo8T7nZQc8J
7Nmsm1iDrh8FvLTso9ut5tG8CMiayyMj8lhD3h23gL9eilQYpeVWnDA8DPcTJfs6
EXUS0RocBmHtHQufoh/HlZdP8Fen7c9XMazXKU4qocx1HmpYHd2XRBtIULzZ0ztd
YLVbk9fkOBcD3GThUKsl/kqE+YsLQ0YWS7e97g69ruWNahtL5MyEAwdektTLiauG
+LHgI3KGWbLJix7F9G4H9ygc1PohtYbpB4KzB0BCv+g4oeiPAkb3xdD/MvA76Io7
nYzNWcGEyZaPMcQBGv+RZM2j+0iTpfZAmMF42iwc7ZbUVzNDk61jj4jP43oTNYcm
LWSq213hFm3S7DMxpx/aT8ITo9rGJceH4M/HrWC9zpMgS/Rr/Jiu2Tg6lKEpPYt1
e/980OkyGVAUGBWKiWi1z6lzPDsHub3kMpc+uL+kh7ULef0QcY8L66CcpOq4pJTG
OBtpWonRY15FWseOMjk8Dv1eDB8ayW/r07Najout3Yhfcx0pcd8n6mPWOkwz1OYs
KmB/hEa+HmJEwpmNX3FjzLTZVM1l8UN+Cu8BhTpRp5R9Sf6krKn5MudLuiEVCS7c
4hzuGTktRTOajw1TEbXHBCLtksxsmzZZOS78NALlWExbrFB1ye1JwWjzqCIw+7Da
W7ptGlUPijrLs2sPNH6JAchMoPD+fx2tumpv93vcztAT5MX2m66Psr7jt5MFXnYV
BrelodN10M+1BKlcnPm/V/ZSlqirId79TTztiNywR3e69H1ltici3n7LDG4Z699k
t7GXtXzfCwwNiZgzuxwGQuZCqd+qTO4Vntpwm57df1khtcXvqUPkv7pUgoNrdQBx
TKvHSIWrNw/GuFH2FoRshTayrsRYO5UQyFWTqiFho4H3RmUuov0nW6XNrJaREcG+
J4sGj+v9votePV11eHlZtVeam9UYsTZhMarHyFntkqA9z77UALbNuci4hkH2YGcS
3YGwhg9047eV7F7QidAhSW7KhFd4Xu4xpPmpOe44fESSP68b05FmIV+g605yhHUe
JHuYPpZzxj7OjbBmF4rk13Tdc7wslekdXyBPthVgAxA1NYPATIBNoDyJIzrP3WEy
fqQUFF+VJrHgN54tqtFqiHRtpnk79H7jJVYmSRnWlEYf+QQm4+XWuM/HBOdxsiH9
WmSW2D2A2WRPLNQN1omXzAtk+4n9QIGmXtT+yVcZpau1wq6PD1q1UW5ByY6ET7ep
TxZ/DMtP0WWlU48slyFyoF4UeLE9XVIv3H3Nr4cnwJeSVCgI8JYWr4gT2QovmSUs
fv0A4GtPAvbYWeybvoRfeujjVqz/9C0rmLVjXc8IfPW9kHFw6kAp91P+9x8kFuF4
7UMGW6pMNK/MfXSeLJpD6NIjkGCIKKmC/B6OFfkOXgDyZF4MHK/yo3cf0tOBxozr
9L4dkBbfOOFhJsq9ATyKj+40b2FiF9jm1Lcok4txyqGgrlD90KVPuxBrf8tpVc1u
BwnufNI27VrozuMasGiMQYAFDgDRD3nooKPvvnVSJpygOqBLsX3m2JRB4LfUTLmQ
+H2BXSHCMY0nW9eCwOd49pSFpeiq26Nnfh2dL96Z4+fWFOUnTInhCZxg+DpwPMEh
rcX2sDyk2IeIz080a8K5j/WxtR8UbJe5euOre5rCkAL8UP2fDPpoB270RlBqRWSL
eeaZvqqGHEaQXS5eA6K1yGQ7guuRlMAH/mzs9fS0MOqJtUFSyjJhVVlZyrCdEltg
JHtfgH/TAweLyYCWygHUTO3FiMbSINyk0xicOoYam+jRhRyFgoV6bKvgzBWnm2kg
ub6XErcUHY6K6Jmd2Bt5o64xmmg4m36jH9V/QZCx+Y1YXVhkOyeeWTF7NrXqIEmv
sl/yiuFlOg5TZKUtiEe42Z6KysOjK0AoJe54+EkgmnkEIcSkLhdcfz0EfDQdjSfT
pe0nKXRBVJ3PsvV1svUb8MZxheIVEc/UVZ9FCyw9VPcHbiVqJKIcBs6fGoGgmB/7
uUS9bYUWlciQB6AeDJ3Qb9jM0j9RyZf+WB0GyA4UM/Mhcfu9ytfrlqgcli9Wv6zA
jnHNo0sDvWnBa070gCxtuuaHGpUj2Gk85TfndVyqm9ZvEVMGMJwLKkCNWcLUBPAn
jYKPkiF585n/phX3o4gfRF338sfH+fIHtwkqrPu+M1M1ARV4Ne5J+ypGIGTkphMO
m5qe8YGdCmiTFS7DbvQvyU7lGezevYsybkdG8HQavi1HIeSFVDsDPaCfaWC787d5
7rW735f5WEQGpP9Xr+wFjreWeDXoPC+JXUxRraytuUE/VQLEaeZQKZf+djp47HEH
T6EqJTFM3UrhkUBZ413+QVg9eklCAebmkq0wJVlObYO+eWX1+qNp5Q7pCQWiESlP
efW6DrH1u5YpaXbn8nC4koJMtfUkfNwife9U/h0STMWAR0SXV0lM6De5T+97iWew
fBxjGW9WcQG8ln2RoT7/3G9f0e69F27kLnbr2SvMCFXqYgWcvbNIVbGNuyWNfBMu
mJk7tZQ3Q7TiFQNghSnTHMublz0lHhwoEyFesPMTa4fXGikzFLj24cqxoJ2ymK89
H24yStKmAFK1dk1heJyXoJMPt/MMWzw55fV/8/oYUhFSVLch2lrht0TanXs7kl7o
YQAv1CMd/9ti1pHhrFGmKWDJ5MTopv56Ahp/j3hk3iVb09Z9qoNsoRujUD++oR4B
81jM+JbkNWRQ1CCPMTVF8fztgpORa10ud799+OVaLnao0MPQwN7AH+ZH+ppNPE7I
bIk7mzaG0Z+HpPM2/aedi15AZX4EOHp+rKizUUZzZdYV1DS1kKNVAF3xK9eAxn6b
+2vClHjipBhyUuwlSqTQ/Qr4uiHtUzqWknZesMP5RrvdlGKAP2DLN0o/Dtc0HK1i
RT84oDtYpqWQ3KHjfHvm8ompLRnuRgBVVqp41kmp2gG0BX+2akyh3THo6uixpxmX
M5CGDKsILB2xqN3buBDPayT/eHxfgl4/IRGK4qJmCE5CxbmRWtLq5Iu6RxxlFXsV
ZFgGftK4pNAcoGzm2tTXrRAopAxkUTeb9CbGKS4TDxDGAPwwHalYDZV/d6SGRSl4
atMx27qyzpb4kliMGbtnVi+GdWW4PDnEJOJCaagTwX1tNj5/6m5BbazNI8t3BT3D
Yll+qM3QUJeQCzAD47VVod4tclfkpD/R9duvmnZH5L4Xu9A1tm4Y7A+t5FUu9dLW
1qOnttRrIjT5aZkbalTy7zHqw11yby10YmfbjKYbuqHeV8pRP9jWcoYdEhLWFK5C
1obLiwyVn+2zxbSd/yIMfrOSsSK/zMK0khxyjIbSONsDZ4sGiMNmh7Ria/Ecf0DN
Cmwj2opnute73JJjY0HIVRdk0IGrIUiOQDM1qjZpHTG3YXgGJxQ4qnX0FdPsjIQo
oujdPcpE/NHCKd/0+PfeV9l98pijVq2zb5SluWWSclndHN2K31dVzarP4Gt6Jc1t
b5QFu6bMXM/ErZMAwtwEGeqx9nuga6vnTdHs/qRJw9v97ozIVnM1ISUC7vRY7ULg
njfofoj+y6KK1ZxTgSc+GB2Ogp2s7phFp4dbdgpEYG8QH2jPB+dAQUEdbiRxxji4
HdpMukaxP6zua2bGcYBX8kPeKgcBcju09WOWVP2QdtMvDgCUTU0GhnSy3vRprm8Y
03lfY9k1VDtmFmKHPQc7kTLLoTLamjHdOEx+Ih5yEerRJFlrqMITNZGD4ukHAvne
4CxugcdDcAp6+IN97arfJEAQOEB+4FIAsPyNl2o1IjfBbZWl1Hz0BoFlZARQ3GlU
oUxN5woaQ7B0E1tzfOcU+B8jiqVtnpW6AC1TyLUBf0JRo1qtgLnyW3ejv71WDiBF
V1toL00T4uuWHAyrt0EbXUxqYTgZa45rAulPE1J41x5o0PWkv80VRTpT6qVkJgg3
6DCqxOqQ9Ss+iKZqz2s3tZkwgCwzeTPWGTJqwlUYWumUmF16cfRq4/NpyfH3F9zS
xn7rSF/uxSmN44qILSKUBSpMj2osdBsm3eJ1l0iNkdqrYpUkVXlB0mXqTwfMJlWx
Obuh/gqoI50kK2kC2TF+MIwBUWq4FdE7kG1VNHVs/+ZV6LUACLcfH9yJ1QifAVqu
LpswQ7TB9XaDUhHV/hHuRAdvxGV53DLxZpn0jDCUHqwCxFY/m1s8YW4gXa7cY/Ys
wTMeo82Oqn9P/0eiCnF42ECWEPru3sZ+47Is3Y6+yVREGFvkF+7Sf3pUF4btILGE
6lTmRtiAy/otFPpyoXXU+mR7KXtnpiNMnu+MHSxgus08jwF8pH0ZWO/RjSXEDhhk
sLWlhWh0XfxLPGN4KI0SdF+5uTxoig0wxFsvrLdDvmyGr32hKqgIPlH8Wg17Ikox
D3Aemj4BAczGtd/5y1NUwjamd8IO3HKmJhhXB9MAv4xMIj293v7NrhllVBeIJN3Y
TdwFMKIG6VxYMW+r5v01nG/zhQqgyQRSnVzXI63ATZ9yEqclzxeHSU2UQb0ChZb6
qNrjPjJX3Hf8TJ8uhyiMCIUO/PU8pVESq5rmfNp/W2fh2jctR2eD2CANHQyNhC/4
j+C9nhYQD6c4T2gHt/pWK+TZf51ekX5Tnv4AeunN1ISn75JhbL4UdMBsupd1mlBd
VDhVpemCrXyrXt35fiJDqlCNlEfSvXtfxQoYoYPbQ3tFCy6SgM5VLiZzMDkJzBEm
06OrneWWC4FIpty0EtUX6kpcmwhttbtQEms0fA7yQX3OVMhEn8F/kAf3nWl3+OHK
Z7NYuvN/TDkRW98Mjk41nv0cpRek4rBvtQnNL6dI8Eg7yCZOxMtIrxKdXL45EBEH
CkfUM8oJkUduL6FbX6M59cH8UJuzQeRRQFO6ktVbduFusGP5eRaeh1txbkTRGl79
r7ynVagMZQ7QLmOtY7zD+/wLUF1njAYXhPdHyOaJoMpnmpW/Q8F4sFMLI2hH4dRR
0gdaDTW8aKQEhuE9UAYYs50LIcAi4LEMpWfd0jMfhaDCutzaxB4v5tqttNmWRMNx
+9boj0QkE7XowIQOEJHXWc9CJf2924G1ww87EsNwshEaxfvMlHykmI7yHKlr37WS
flEPWAj6lT3hDQaldtjOknMn4dbDDEnyJOZPm/W9bTe9S+d0OUikgU3y57NlvGxI
tYbTtxnZoOQyxwdjUZjGYmV/nE1AaLZ4AnZXdcNhxXhRFsNcp9dKAFck6t8Ia/ap
bhI23JAdgDpW6YST/jxpaXn6hZ9TX77d/KykKLjBDuNnbGIQ1G2O3pDyxMzGh6wu
2qkZnmyEXTA+a5tWkpGZWnNWDehhBDxPDZGkKjRZdVbam0XCcULfh1Qu0vnNGXrY
HBJbydTCUz9lfm8MLp/zfkw1Q/CaQqenDK2b7ROjPTo7zxg0BDVP1fzyj7dQRX5H
W+bUs27+p6x5T9PR98uRqXBclAs60/w07axNI/su0uxm8goKnyRaXYt9dG/NNBcC
2GQL5UgLwhYrPtTqnqtfKLI7PZwrSBTtjn2ipBiSZP9mOmJW4NbXYdzx9HUIXjrg
s4VlN4qbPo2wFhUpx3ZYA4uK33agSBldo8WgpTXTPmP3qctHfCk1OyZ57p9A2v0c
i//Dc6KKLXWmiFnEjhdxr9LMqLZbaLg/zs7rvc8TVrlAYtvkNhep5eieVcv0ZlBH
hF2W6/hhOjfJvKReSQNTVfTtDlrMaRFcG8uZ4H5WFcP0cuGWB8yALOccMzoyxXKL
Jju+LW4uFhcDGtkBShDhA3G/An3+MQ8mVtD36ZsJmsGebUglO3pTmc+f7UPDXQ/N
GOJUFPteiHk0uZea6CZkd8ENrPAQLs70+vqNhc8aygQ7qNJ+tSpBBsX96zg1gd75
mwdRFrlpqI7jSjYBVYnGvUhG/sliT4ORrGANZM4rbAYPkpuaaEA44Wu90eextL/F
GbmWUEl5ikmvYyYcsc7ctFXgksTeZ4/JbroVtv3LRGsGxP0JmcSGVEe2zZOshYo4
6q3vgnc6jLujSkydRkMZsiORLVal/K2RULZF8fn9MGTin1QXQYeHs0cs5mdx8JjY
aOqOKMFSB/ghP28qANt425A/CEFBq3O8xHD2GTzJK/g1yPBOgFxjgYIp7buzYqYy
Yy36zc6YdxVtZ5LVsA4tSimb36ion/gQAxY2sSuZPyv7fINyjIgPHuryMei5kXol
CDwAqpFZTmJXZJBE88JSMaq65UoL2uy/5DJiYylxnWPbYVBhpLZ1LPFglqNEpTYO
92a7jnIGTvw5kdrJZG/8gYn16pJ3fggUUKdaAta58S1Qr3pAUKr4Y+ZzLL5FT4Gi
TyxKT8SHHBvrWYgiGa4FYqj/TjPYwbJzmAP1GQPfPJIOu735mIFft94MYn9RNJMh
IUu2XX5GkPJphM9W/VbCyDCXD0Ziyyu2+tYegJXLBIzZVAJCeeozuRy6NPIdVqSl
BPcCFn6EHa+O2Q7ygXCFxdBTvArQPJXZxUxIwjeaa81STfpVFhATYu0S1UTnYPq9
ZIreqFUQxhCRztm2gfRm8D7eei11LwL6zvqgfSL4E4x/Gz+P5qpXQAOX7Y0AVKrv
25zTXXTvVE6iYFRxuT56ikUckUGyI/js83a5yrC0lmyVeWXeLLJsZo41xmvZ8hN0
uXqZFW+30sk5Z6QMzu5595+nDonL58I9lpkL2sBD7iiNj6R0pEJ6V6nu+pQU4/1f
MiwhodqcgBQciascZhO0YqSTWT/946wM7Rp1OReSF03wO9Abs2v4a00eh9UtSpCI
7edd4Pb2PyBpq2G8t/uyjQWcXemsNXHOZNJGQLozNPIK7i1olx8yerFVp6gr+1Kd
/BAPvNO7dR7wsr9SjmOCFkIkIBVNOi82a+ptFQTmNzUy2cnvvsfgR50l+44BC5vo
QoHGVOfLkbGDZtC45wCLbVLXNjg+zpcHxl9gmchh/Fv/G4kjZvezCbyVzEgNZedh
rMerYs6c+hliCKwV8E2mmoKcXwBV4/t53m8InOhAWgSFtnaokYriqz4MauD0vHA5
ktHmnzqk9YoEsJ0e3djyYVTLtNvzJB0a+Vu3Ih3At0wxxmv83uAr3n4fUvZCdpL/
XCTMDjVxGuCbUh8Rm/eNpZv1Zlf2rXiAcZl7USSLsOWdCnhz+hJOLhFSAaxBVlyV
+KjLe+yViKVpeg7KJhH/xDQAkHBchkEaCa4ObZluu841tTfWBOK3e/1L43M82dQE
rRHtx+svXPDVqNaPy0FcJgU+fPlQI9/HRwwSEzF8ZxD16f6HNCa2zKFhnIH/+XKE
d5urV/saa1u1gsxLdPNYB2tOJ8KAmMUruGNlFcRSVE/JVtbp5qiVLVFyfiB2HNG7
dmz9SZFOMwvuOXMJI73Ex5YKCYsvycH2G5Dufsl4CVxbsOju/oLWKRZQxXLVC56B
7WyEVuvh4WL+IF2EnPs0G/UD2SZugI5RVgILNcwkv1rS2L36GGZ0+ULuykfyQV8L
JzFVdliQSk0UU6SZOdMQuymho657gpSPj90a6R33Vmqj0sKnHql7RQIGSs36KHDB
vaLP+45hCXCj3TUJojii/Ys+Vbkdeii8w4NI8Z2A30AekHubwZv78nxV1CbEy9dO
kqFufpSO2A+rVejKJuJYSsNxIe1bEJj1ZPOrLVVrEWlqKgSYa4tVbpgKmhLe8zZy
oalbC9rocKIu/Hn/25iXv1XnzF7EyLY5ZvSY4/9JOn1qwE7xiFwBTmx44xyOU93X
GIp0FzImStns1ySebOeI1QYlB6oL0RCpti6LVER+ztsrrtuRllVCcmh0UyTrOsys
mktCaE1XT+lA5N+StdtvvVhHZatM2liLIRLo/UQPwY7pDkntRoc7F0vQHxA3SB8W
n+qk6ujV/068fP279CNn4Kf9jJ322h9eZ8IzdmL3+cU5fAQA2OBWVhbBeKk9cEXv
x3MiLjsQfzOVPUTij+9/r7pXTh29JU7YGFjsRg7f6sQ4zbjy3BpE9FwBrPlOzuxT
A3zipExmFCFsYhbyTiq3zHE7nNIY+wFHfao/CDDqzlV8imEsmxEN48VE2UV8BcKr
uPqmLfmCPO+GZXXpYStCII4nh8evgftQE9majQl7ztT7V8wld1oZDzv8ithuGyCf
PwgazhtHF2FcmHqaclEsAQZ8gsB7autR282yg9vxn715/m61Jd+xhp+yRlEhXFOR
vVdVWSw4Ad+06eLuchBGich5SwgzZijcqZk4xmE7TG0GOcrlISxDR26Y+PSHTkeA
wS9Y/21e/oaaQs4Sqo2beAaF3MEJi+Y+M2SW9tEXUEnma2OXTZQRvRB3wiYkBCKe
88JR+cV5/1yc5xLeLeA2mgLKz+EivPIhx9ITdHO/L3wNk3V9zPBL6fSuUPgL8Vyz
7r42J8+CRJEvkQZy6Flf88xJYuvJj9Ev9h5l8cCzlJDaFjN0pQw46POUoqip6Oag
gCAumgZJfjSB8beitLEaxFROM4fMuuCIwCbXMJpXWd6Azh1X7eyOKe5HxagLyXEA
Hbjkl83qfNpeWsymVAs45/wWPKMjlgyR21s/4c89woLUsrIxmFPPD/JOGpQvLKBA
wAmDd86ybekIMozAY13SwyKT0gGD8BurSF4qboaabNXq3fVj3rloVbmC9NZZdFsz
BheFHPlus93mv4jT5HwvdLOD2fDngaIBdzPLyJ7y3xB9BeEqaTykYxQgtfdlD1lN
sCaRJaW2n4Yt8Ri9peFcMt8/7x0RshjTI4eHMxWe3p6R18hKEJXTE+5L/WCaVtOk
SNBTJZ3ZoODNjC5wNUmXuRWxCF45NfHJo2g22nZrFWMCbcFv6r/yWafXraOR0vZi
B9M8vyiuNIJWLEbZPU+8LWTXgYACAvTwAjUAggObQIBvs2CuFA72n9KlJzpLQ5WX
1vUqkiutJwKs+/d9DJnSdNQdmSz44yNuTIQR6kbQ3ERGZs7wfp3OA2dOn0hCcoFv
vphHOoD+lI3xPyNCAXB9FzqVmzyqJ1//I+jBhzjhqvopEiAdfHl/rU1hghp9Nd23
3uZF3wTLflHFNwtpIMdilLeHfmGZX6xPd+WqzPH9yuaDPL6Jl7itHvymV1iZUgH4
+lJbt7P+gDXnWZD+QgLRtPJb/A1y7JdWeqbLBYbud13LqCc6JZPu344Oh1Sl64H0
DI4GfhZpSApB3a2oXFXaJzqjNwgk8QmzAxkabB15alhiN/TqSX6dTzNnFW+xAspe
ILTNalxSuW6W2TnwQT0vEQpjKCo4NTiRT5Q0HIoTKHMGpNkHfc7R9ygzTp0woDig
9dAx12JZTjS2MPk2a7oxbjDm9fR0h5bVO8kcKtTiK7mVoXTDU0hba+ATcO3Qap8P
ato2PfXqb41CO3SArJuOYsxdxV45VTk/JgiXblWfksJcXhdNyYOlzs32+8mf6vj/
cBksIMLpM+RxUYdt2ykzSPquvas5+snGcHP2RoB6xK7eAIWA+doIqUqORKhzRrx0
suQxxEJ/iCjAyxDzfoveyHBMslpFtY+lJA4AZlJk7V9EmAFvr0ppi0BrrvOqRSBG
oFMziVeMN5NuttVrB6FJ+qeuGYnesGm5FT7JS2yhBmk3ThjBa8agBk86hhGAxseK
v+JwRuXNX4/M1/IBsZ2xRT5e2QVZKcSAFWMz90mX5NPdPLmnLgr+AA/MaN6TzCw7
4SSrqCT/FHA8fCfRWqijSz6YyhduUeuPL5cZ60l4mtYSGI+WrpDHNERWnaT66PeL
dsNIhnvGnHLhgl7pGHbJ4OghLfnf+/IIAjMF4sPCvMq3z/BXBe6Sm8hN7AhEoHur
AfJ5a9Tha5o61ZpPQYgYYj4YIN/meKFfCLLgWnNtWRz2/ib5hVjEXutFcwjKKVXv
oWAdpCrpdppemQLdgjW+Q/EUVU6W1vLKCTBRZRs1VTqIr/y1m3W7yew+vDURkytp
e0UUG7PYEMnCkHEHi6BPtVK+MKTdt/oEmGuyc2F7FzuufCmVfE6vsiZrYgegyX+6
qZouU5bVtp+hQmIYK//Ei/uXb7xUDfrREfDkV2ubjz+vemASrK+ucjEGWoOwSmWW
MSfn5+r2DMZ1htFnWqq/zno3aTXSfXzfUeB1rGm9YSHsQbIEsGyxv3bdEOo5z4Qn
WA5tPxkaEjor/6vrs2g/UdepBEQdki6lrha0y3PUvBVhW87v8i5t87WPgjr8oigO
NonacEF24lLpaoRrj1vz8HEsRL5JpTySwXKVnRg8k7APzkMoK6L4KWGvCaZ6p0Tk
AivxV6hipX1AHBjH669etOz/4hx3jDLA2je38M3LFDHeGFLN5AXBlId+XG8evAZJ
ifduan80jpjg/hgn2RLcOrZ9T+xtuTj2pErb0eE73Q1P2XEXqDoODKQBCTtBS9Uu
A/8N2o5soBjfST7xgYfPzeOcN9SeHrVAYGRqpTkFvwyFG4HSjJom0eautIovsQS4
hKAAJmauPryiKPIQBFj5kWc/nwbWy7Xh+sLuSQSk8uvY4Ry+CqV2RjwKsOKNuPob
YGBzk/eRbJ9fOd8r5yq2SlvkIPsnytxOCQBNmR/MMLh0Ut4LN2a2pXMRHV8MwtUl
Wt0WPoQ/pb+knrAv46BgGw2jaLcrwUwIseLo/WN4CW25/eStA8wxRH5yYd9YiKHm
mYQTPoFXwrur3jK1vuu2mK59HKyHDGYuTtVeqfaK4sCDn89zieqCtCSiPiDL+1qZ
JD/6yQHfTyKsNc4TlmNQfAMnsumOya16lgolgwiNaV6HJ48LVbdnivcPqQfaRedS
fxin0YugrZ3zYe3i65DevZ+tEcKjcCbChGTKTSiwypVJTTWRmL0M7lkhWXGLrbIG
Q0yedEYmx8hAErrQZNTq/nqJoI/8E9q8xYVxlSxFNCbMp5siV5tkCZwT31Y3IXD1
vaRjQoPQPCE+Sirmji33iJj+/yDUrlzKJvWTVm1dxZ9rCGqBqIPVJyYB/5DKwmEu
ZfRDEMOaKi1vLsul50oLZNu6hQDf5ju/YXgJ1yvF1mK4NwB33OorrIFdQJYOPdGC
MlZsKYUnLMYpmlHRr5V49vZY4IrDWcyclZK1BeF9u+0ckC3X319drDYA0ri1qhR0
Spun1LYU0Yn/E52II2mPi7p8N2fqCvvXDyvU/WKjBhk2SBrC4Mbc7KuioMVk0fA3
+aIwJU97WmhZjuCeoXpMg2EiRbTjhFkN28u+4b52TlSWpH0Pr2C17kStm+Oeo0Ft
sYaU/xg53f84z8mXTgBLIYrt2P9dzVmE/eksBVF/pjl8tF1XUifGwY002DIv/zeG
WHb/bHVG/hzorK/NXcT8y7cXCSfq/ZsHaPOWpU4dxr7Dz6uhuagRx46bPIz09xdY
f+VguMjJQHce8Kb8PCNinZQTFBoL4xqybF0ntvAwBB4y2psm3iWfd1tzABFr5zTG
XlecAdvBCWtszYZ8FCn+HBc/Jk5mFHPByPXsWSi/jKbU4KIeRnVGa2Ki2HLPPqxX
HgIB6D6vkwcx+RCURpUCkO8U9pLAwdZClA+1Z7xyZWp5amZBzkMIabXY6qFAUoPa
3yy9+QbBv8YInhHkEj8wYhG2ax6h2KiO3st7ATyUQ3J0PhZ0Y0hn0B5aB3ocJFLL
mqAqQj3EUPT1dQ7v4UrVooZZWdj6Ggp6VdZK8OJwylYbAPrWidMV6e0SQRdPxa6G
GRG3yzL5hIaeFxJl8h+0WaYeZUZQpIDBoZY0jGA2qZm/NJobawy3555Kbu7QdYHv
o4ikV1rtqRUiPgZ1avXbF2oj7FJO5FTs4eulzIq9xr7CsrTMuZQwCF+Q/qw5bQ3v
dn2qaP41D6ACdC3PMJbnUuCAjNQrxVZmPfu8BYRn2vvYagSgEosQv+j/peJu6TTQ
HGdY/hUEGhs0iaS3b50oSfrXKaoMDTNCat8fv5yhKBLsrG2HqjxDuZkarRxSpt/1
VBJ16zqukMX/DnkUFVSSO8nNs6xSlJnBLEgPJ5y2fO8LtUD7KiDhXsbDydjrirEB
RcsRcxWUxo2z2knqq/UWHDXsCb7cQ9Bm36GQnItTWGPrCJfq49N6SqXHAszRZ3jZ
0UKdrN9374qeQUnV2YUTuYGWNQX2rY/POctgEuq9i7xMFHT0radxuPYy7YNYmC0g
aGQhMO01wQh+v64p/1CK0qXfEjfRJOOK+zt/EHH2n67JV5sBhC21mg/PFBzqneIZ
MJgXKTnvk6JyKLlX/CJ0oUktuqdHKmKxaXI5tfAfA+hEDu0/TeuOuZl00ZYaxlSX
l3Qdh6Ei6lyWFWH+MuL5WFAaojJlgkz/GWg+gJ4ojyp2ozU0v/kImLf5xnEHW30F
p9d7JCu8jkhBG7effQoRFCGVFwVdplBih8h6H6Qpl4W2+Kw35eoEz4I9uVtvtwLM
cVEGw8MidKdLHBO1XvO16b9EEW851yJDpMRM5uDZVqMUYlAs+LlpMXYNUodJao0U
CeOsCdY1zRWCjMvJYZC3Q9Kbjh8+ryhDPQSc4jpvZDAJ7s3+ZFvo+utBZ5Ule8Yq
JEc4kVHSs2X7mhkGUYCFSbkjYUY4b5HXiBq4GraWhCrAB46tjtiea3ikSADA+GIv
L+KHo3urgRlWe0usFg9zj4beaQYx3r2V7eIRNedqyYNeknrE3qX8xF6coWDiQjDC
JbwlSYq2LsO+qCkAsj6WUIs0gRE4g+I992ua3dQTD7i03PZZsAYh+OJl/WmamhFL
7yEmdcEYx1khuPaIMPrP+Yc5ZgMpOLmYEs4eG5Yly+6gw0cBhjYQ+AtOb+DQLKxH
Do417yyKcqCXHEN/Wp2eLyevu/qXb85Hrzefvqzk4JWIEzyND6sQcCZPNg2jHEIF
9Uti5UZ2B8/BRDil5uXqHWfY6hiJ0+XtIq5zpCh1qR8t/zr1VMYZlAC2lewjW+lW
bHAzRQyqMYwK4JVL0MMz7iNnYt2mFUJBkRfFR3lC/okDVJFjrf7RD/pcJCP1828e
8JXqMu0cXKwXqp5ST0TVdyrplGd5j4p3itQ4fX6N3qMdkLV59IOaHSAENPbtboJ7
WwS9jkRwbQ2D0aYbHsIEzQb9wHpl9cn14kp9BRmdDoe9IgC8+KtbsdoMH3yr3Gtx
xVxeqHvKJNUWwREcHy/melt4qaZ+XlMZ0IFa07K/GW1kkPXaU57rpxvlLZiA2jlD
iG8z495efnpYr6700wJarNU3qQ3xffiW80p5/WZ7kJiftPo2czmvCeE2H5iKzRN+
Hmu8M/GR6R6jHgXmKA93QGb48NNepg6SpZoMjxSOIKyiT/Q/bwme2hvJvvEU4drC
4pQDFr7LaA6fZ0cRq1ypk0wqIjFntul3QhWbHGP2qC6+glZQAeSSpj1huHyhn0Tk
nnj62wvJkLOVX0EoMzHauWUyCMdcg5XESvs39rkSmRAeRJmZu17Jerb7sAMItomk
c8kxtjrivMBZpmJ2p7MdbvRvlxaJO+oI9F6yWuuCvcTCDTvt9Bk/0xDf2RPemt8r
4E8ZaIDhjvyC/r4PEhA/c/fkj2AnRGhufNZ2hDUczr2gU+pV0rzH70wwvraCpgAo
Sc6LpA1GuNpovugNi6D0IyAv/DJst6SEIF4IozRegHBudQPpq0FB38inLx+UxNvJ
PGKt3iW47RBjJu/1Rj0uUmqRVvZfSYXC62+7AIXBI6OZrgUJklczfffP2a4AsbXl
Ed+bwrObM+A9EQqujInp0DVR6SpuUbtmKDQne6n/ThJNc+DhfouuKl/8UcrV9XXw
UazpZ06LBOf/bNC731g+52YEFMhYmS5EIr5Al0vT7CcftNLJ2F6PZyCW8J3Yh8Iv
nQs3XSEO7RaIPwdap0xk4tqbupDYBG3YAK06s+Wp/2QqJ44X80CqORUcYW7LA50M
M4pjDFAv0Yq3zcgG5tdlroz9lN9A1dN0Ysx1wy9QFqG5ZX0rYzR0LwcD+JTJilx2
tEmScOsZIVCBtZiQtryaRo1LsObGY6ZNe7LpvbpssCk1jgkIGzMiRPgMuvHRmDn0
JkRsSpwrzdyqqtykrz2fgNl8kpGMua9os1sdO1EkFLrS+RgyaCkKmgV44eLHBIlT
w6qPAO5pikuASVQeuH6nafnIAP87y47xg82s0mUFx6A/o60rJq7cZDDwdsPLn5nv
XWvE0iNXDynJqD+LM6f/bw2yVVqyxJnuzpyiFtPWdVmIKyBTkGBjS5KCxt05Kdz/
0dw5eYtB/E6gaAA+WwJLH4wRTSg9PIf1wFGaIWC6CCnoVIiXGGPsBoDNj4sljZ7V
w4K0Llr6Fr+HZA7DPEBGzHuCUyUk3lQlgI2ZF1T8Uj+AwrZpRyU6JvR13seKwc1w
lKQB+NdVbb8GtUBp8RviAgFJhXBdedwuMvxpNPiLHwwrFfcI/Ig/pyjiKDhBJI8M
YRPZlSNaGGPd1J/VDOFqeqNHRXgmQ7dhpEBQByouPEcnO7EqH7buwWaOz5Ec9fqU
t7JHO/DJIt1nK73X5/fowkEq6pF+xufuQ0WFFzPx/6yFlkP7bA5pGtxeVSsedxo+
gQEFlkdVVzk8bZciFH6nXwnFn3iczlNcs2hyfcvhu0ThYK5vzt6X8UFVl0QlhtZG
aybSANY67PpdQWLMesFALpNPs0yUrwf0L+lQySis3Ikkdk06BKpUvw8goEmFroq2
LGOgKek9LkCGkPpYIxXHNgS6rx9p1IxWaSRf1yM71Q8sUgmJxsVj0Z4U8rQwTttS
uU8swzlDiJ0VRN4L6ZYNvkpnOqNqspwLU7tE4JyzLMxlhqt1Gzi586VVLEmW1Scm
nJGaQpBWB/c54z23vvoU2hXgDdpy4h2e9I/QA7twdDE4XdeIobr9Ne7vx07B/AO9
N4zmtvCEf8jaVaPHpQpxH1a2M97MBg107G2pWP2uV5vE++zq4yS9oHdA2OmouBGU
3duvPZ42E5RH7Kk7YHp4TMilf4gHhJIarOXX9vQSKA1dKQdTbNCa6RoT7QQuqvK5
HMmdA2Veg6iKgOZf+PDndFM8ENGuGOoW/n9uhTHd21VnowclTiFFEyQ8QgiHOXqO
rFkUrnGOpNNtob6e+iJvK9ZmJHi3tZUgf9B7bO2RYad0EjYi8joXbpyhruxpKAV9
eWHRy1dBqch4vbAOBNKzdGvmYTv+zSWwBLMFlyA3f4rYA14hGIZm9noDDjhh108c
WJi1OhsSfEKgBS3WFjl+vwMq86yh92j1XdgmN95ekJ8oEOzCs7JIZffvNFdIRnsX
1Wk7JOPX2ewOGEHPl3GKXS+qNdDP7rK3bpSP8KrPjk+qJBekhDRzf/UZvNuUhthm
6/ONvYwPIB/juLoDEdf8tUicSy1vF8o8GdCe2tM8nNKR9D7tSDljgukVvlX8gGzY
iMRDR+KT3BMJjqhCiCcoNkMYk0+PSliJ519G6WQ7ih0nAOYyTU2bFy2G9iYUDVKp
MvSW7X8VE1yJox1vPcPy69ks/7FJHjQFaTV+1uJH3GiHD18QdKhOwdemWtTz9zPC
Vn+Oqn/VRwmhzU16CilvsIo71A1ELkMriD2dCpQE2tGyebKGFTVOYeSwEWSuiH/2
0Rv2tkGl2Ho7yaswH78oVRUY0MV9BDx14dHOtKIlNpUk+bo3sE9WPEbKNILSQhfg
+yO+1Wmc+2oCBYg+bRuZFHW7jstaHY9Or1BWgJysaP7RMsTUDt4x+3WrD3/P0mbX
e0Pr1JVU033OoYBV2JEXT78j3UzyMIbyuOh/SSV0DILPO0JXWEUxbNFspicI7tsC
uU4U7GgIv2D8c1ytzqTMZW0cXJ3g8DcfRJH2/QzDw6h108g962jxlbaI9nDa/q/H
PWb1t5i/icXkkFvfEepo4VidB9zxnGSUYPb9jq7JM4jXiKYtGVS4U+QWq044OFCY
h6FS7706h4071nhGBpdAMpABC0SOjTRBCsVKD87gWdOkXLq/1toQuhe/5+kY5XXj
ZFLTi9i54UKLtzRUmQYjzX/yYgR19jD3pjRyBNLDcGh8bX3ACrz5yHZZ62DUDeIa
r/BIhsFUfLekmLwbSqeOLtaimwOvcCUF/8WTscWdI+rF9qKszFRPyXDPT8TrAvpI
NVWMZBR3bI1aglKm4p4v8kRpgSTcVBkMoCfWOUtfLAn4XdNN5WZDpTtPaD2Gh+9d
xICqogSPurI+UjLnapJaFmS7DZTNJrB9Osdz30agGLZwGr4srhS9GWUHVPheEXxT
EApuWQKQZ44eBqXHd1b04IVxHzkIE0mUO6Bh/AHl568DeJZmTWDeNLuDwdp/ZoFX
JsjmnLguEvG5jRmePRgYaXIWnizLXA4eddVOBRu2qb1iV8k/Vs1+wRd8nYElmTla
DratlOlsllJ0vx8lTIiYIV2jtVXtwd/ohGkkhCRp8+9PhuiIAzgcY+viwV3eG6Hc
2mXfTSzzN8wL0Xg3e6/GK87k6KZykBFUKpZQ6Nul0XxYvo8t08XC6FfojdSblbn7
mtHSHb665+bmkoA6cz7oSqdOr6gmlknWid2kwnYAMYd7I1yIIjQqGKk4Wp6CmDr1
r1oeB34FMpsIRUJNUw4hxICb2ZjXep8sUWeMwxM59x7HBm8Uus2VdUPDD08UKKuY
YGbQ54YhsWKDi6epe1GU3KEwUyNabOJ5aod3npylK7raB7QcIXVDW0dqMr/4IfZI
jLxa41mIZ3YYho4gkMHjBXbWc+j9/9H78vTXUkkQd5vxdmqmXPdkVaWdsxiVvl5I
fMuncZl91E2ip5ScfxwzZSMhzN8hBN4jEUOOh19QdGohFbsJLy9EBhEJFW3feffk
bG95SORrWnjmzXLkL4Ey0PafNcJ70kc8StloULa9+uR+QN2FvWf7gVAlsyl2IIGV
PGx8Pd6ZL1jxioe4irZGXOkXz3vKyEiHxLsCGivb33SPnyNiSwi4OBX8FZt5k9rV
SIdrwFx3jpYwUNU0fUCwse+HX87F5kPo5hKFBI0JLAwhbaRfcKv15BZJhC+SMXrD
TZqVPnxBhOQgHsSR5r6YseonxCgmdsXPiVqiZdZ/9GUBVKMzvYlAc5K1wD5kWj++
457KAyT0mI4VnydIRgUOB2xvi1PDcQtYciiuDEeA4OrHqm+eKOc4lZZCLpY8FPCa
i+fQ4eRGZ6HUILS2Y5hjZyGVIMU5k2ORj6nyGVBhYFbUHIuJKthaHiYYriI2/UE3
9EbaET70M3oKW40gw4sBO2paqx7ej9fBAj8NGn4CDKU/A0ZQc1r87bH2RrXLzLPi
1Wnuik0kbmWFqM4bYhTT3wLltJCyx34HBy5ifPYDlbGhUzuyOd9ldUbqWTIRfxmb
uJ/bZZPKMtwI+di9FSPQvAmufif3u4ZGPKGiQpw2542mtuTIVCP/7aBOVmhsZADX
0JwEn+56jvoNyFyMaLHo88lRxxvSJIom8alE5l1SFcHdq0Uv7eIjdww3FuCsOIDm
AHvjWr5I8/Ab0641rdPhCVyQADCaxCtaPT7qbWehJAFHXUlVVd2ZOYTFQSLcIbzr
nWEWR1EIXao+fhANDIPTZCGAiCvRwy+a9bshIsD8H28SCFeqkZtfy53zV3dX9t6u
eddorN7Jj8r+V6W5X1kxtaOWAyHiBCWg7Rk0F3T4KxF62RB2Ham4E9aZG4ikixcr
m1ThxVj3yihGrWi4wJKmdZ/RcNC9zcMW3x9AnJVwZFoo+FC9KjJtmGuoITcpVNYc
pDH4qMRLLCKE4K6dt7yDPV/r0+NIHVvN8lGo/zKzOlN6M5NPviXA3txOnI/fxMCb
+pF7G57NQlQw0h5fFjVuHANqbGXeyuh0w56byH8TBvbp3jqBSCsuBNzW40GSDSyB
7288HC1lHIBZD3Su26h201sHReZwTNdN3piERCFsfYa7vGuJ64zERrE2qypGBrmr
RV9W6R/rDyifi6cJBTRE5+vG1bjCoklaOuSllrLqT8KFFmzggnX40KCVLREdAATP
MmgbBBlyCzODL0xMeIL+M0EfN/cD+HWlOsucC4RVerMGQAqSIGJQ1Y+sSpg0WHmF
iWUrFdwsatZfl9FR0K5oZ7EGcECN54utrRKcSGd3UVLLe4IpIKzF9WSxgWwa3N2b
muysHyYfYQxTBJ74tnspBN0IBKioGDnEnFecVZ3mjH7c1MHdOu+U6t4zzE+JY7sr
Zti+q5zcP0oZUymzHEKPAi1TOoWKw/jycuDVOIrER3AzavtzKPmkGKX7/KnFBD56
7Ah3qFt3KmfDT+M0XfR8vOL11hmmP/fmJtwcPwKxe+/SQE7gLPXifFa0oQNk/Nq0
Jt+wT9igHFDhIi35l8csyrcAAj2VgDtQr7HHky+bi6nQN7AJXkFJhyef91JSi9Ad
i0HTlSxncpIdLr4S2UCS6ND1mNpP9G/ZpOKi6a1VwlwFog2kC4qdOiGNktxjrfwc
ZSKiaeGIw6z2pSGK88+pFZO7oQ2JEV27LBSJxENQUzRzv8ZKY2FQz7Kn3FwWipWb
YfXQRtolR7kgGPrH185kqn0N00Vy9WZeqWeKIgGuH837/k5rqX+A1lK77F9t5f+4
C2B2lCi2dVUOd4RSlItIVx5b6ihHjUzvXNDkzIwaz/E/c69i0oU/sksKIfNNuukn
Gl/oF4XzWGMcVJqKfWL8/tXxaHDcAXcCFGEnFSVPvF5ErEuCOLvLAFuLuumV9GMR
z/aEf+C/sVhhXc4pERbnrot6gpol9hZHJkkzMBVMBoLFuFsx0v0er2DUfAkWZCND
3O5jhofltFZ/kdGsl3wo6B7M0J0EX1hvwshIQmsBgSkBAbyfbeMptqnBV6y4MQC4
bug75XAbXf0Q8BZ+O6NLYcAFr/sef/MeWE5rys5u/7eOx7pYzTNpLCKBYYfbygxz
kbPlqfKTSE6Bl+M0Sue3YbB/D9j5u0ZiwadcDV/WdKVNFFJ7CFK3iqvaIvCfynxz
j3rBLwXTuJFNFQIsUxgSCcUFulrbL0CINGA5NEO4T8tdukXGg7h/s+kpvVkfsQVD
tNd2tU8n9zsoEA+1C/mIodaAx8PSWUnhyzbudlJHb8EQM92qXhZJ62NcRW75VFt8
fdjF/Zb0E8MFayUnrgS4NjuXNtT1h/ermkn3q7OCqGzh95lVl9I9yUKerN2jMK3K
25d9VCAc8E9qXgMcD+5v5UmXArjNiDw1UYCmhIw7a+vOSXMTksY8mCTeWUOSXJnw
1iR2ZLbGwkRZC91GAuDdDPaO+yCJCuALj0uLkcSgX0aojaZOMC3BSpeWIe00cakJ
7yFcK2XI98J53UVTW0RFkAv2iqr/yGPZAOEe9QflUMLELqnCJs+VbSjSya1MZZlz
MHIzCeuQ4j1pBNY3nLfyHh1D0rBtLqTBzGEtD5DtnqvgUWe1ibxA0oNUZvpsB9wJ
iCdysCQZLiFjTOdYdFlalRos5CLBHfRmIbFgsMID71LZNUcFxi1wC5Th1DC2i7bN
SeqCpvu4PWqsxREvsUHj7JVbWaNED7QbRN0C9ti99zm/7Pv3Rk+pYVeBmsnKFT9P
XOSgW1IlTnBNq00XnWTludURQXSpY3lLmwNutfIfbwc5oCC+GsXE1NAtCyDqbRGN
SFuBWEs/TChBYAh2SpvsFYDgC6P9WFIGY0aniD1cDO5nJ7w3Mw1E6gnk8TwYWA7d
t7cd+N2jNl/EQT9W2aLJIJL4YmVHGxNzan34SM16klVTLZS3BC9MI1+uZFx6YCDH
voIZC3Dtot2pOKBE4/aogws4xKJIHbc9K2QLB7tgj4rAeQ0URutHWibtLcIOhBSh
nG/cHeOyZjvrsirsL42drC2+U930ROpaOtnQJ4r6NAC301C6cbP3Lu2P7NJfdwPW
vvcfSnXoixHX8Yj4lgc5aE5TV+7wAxNG910tbYoLjiJFbZQwfZTXmzXIP/r3OKEH
BOyrTjjeNjk8xVq1HkgzZULmw4e1MUEV4bgdZBbV0cUr3SuoJsVknfLmkoyN1scJ
dZBZZtDGT+tQunXeUvHUQcPQSQpLxN3H9F4ptifAfpLdDetFH3ACVMOlqyJO0vki
qRss3VRGc9xDJi4DpzpUw8kW6DyZzzZ4L0kgLrFky18qCTCXg9tUYpqHHwpiqlWE
q+ucNOl9QH1CBZEbIDB0hxkxv5c/3ajbzmHlc2uq9fQ0eY/vcOwcfRVW0a+18now
czuz+e3hMzw2hTTNQqiDoEKxCTykGzlgxp1yBJToux4dr2ll7GJabqyZK5rglVq2
eN9wsvWB9hKeK//t1OUlqwFTKoD5A7A+MUT07wumlHMqHf+sjgSc9QuFhqUuFc5V
4xqpUVf0tIE6dQgnh6wPFL2d5oT0kvKnwIFbBiC5soY+gj/nGlF+HKzEBdRGq5sJ
T0zgM2uPCpiuZJ6acVaPjDmZGivmIEzLYC9HTqq81s1GwmXAr78NzzxHypITKqie
XjUSWTF9VYB8jm9EZPtGjlIQgiIlDBshfvV1zFIL0T90Ck/kIrni9aHvdIqWmOOk
JDzG/zBfeuo0UoDVoQjku8HgslzmHkVCafzEJuEGFuAgCBkTtqxz7CqAqyZBfE5Y
D1oNxt7h2yyI9niUa8vwlTVjh2Tlr9iKbBB+iGs/HGAdY21rOViPED/qSPqpmW9n
cCjZF9BOfmlNt3sGrAM/HIZ/zHX5Fn5MXJXCs9AeFj4WcOsQG5ITsoRB7lg7RelE
F7fdx1ZzEpLlGoXeCqXW2OoU3S6mwZjwGTq521GoZ5ERAxETr+4AWVvm3Al6lwTw
v9tOwwHl0SjoP3svxS5YJYn8rb+or0esaPGRLlHzb2yb6lxib+SI9XTgfJzu+wHe
rvDedTQ4/wfkcWLIp3xk8TM+jqD+fEPmetDTKg4lnoIadWIBDkaPMBxHdo+yaRRZ
yBdkk1HfhokxvGy0qIma1uvIvNe4EvTq2UEB/IehE54XYuONqlHyjj/Ms3SO/PHx
tHAqHUbzMP7Y759ESXRAzwh9SBKL9JcNZFL9qudt/r85VGgO3pGWYriKt+GQi/DU
+F+zfPGJz9YnQcUcq0TkEfbrwzqLJJdwO6qxc4BulHCEwOtb7sURrpyKF36Gz+NH
W3nksUHhH9wDyuFcNinPAwnmukpnYmGb6T5xpPaAC4BD1YJ4tYclEOcwQEu4OMq7
n4i6vhz3DXOgBBGxouG7pZtAIvXWMrXZk7/kGCgYytTynoVQnqW5ZNXktj7fSbdB
7H/wekVS8fIaJ/ji4NW15nAWh3ed2KwaD4yQxqpJk4AzmjKhRUEFJ8zgaa/WG0J0
ahnaCoFCId03lbfeBFd60GGpCfrsp16t5t/nQj90CM1JngBpVyO9MDefx1uQSBWs
c2puTNhJV4y8kNJ0dnriOCTOoLslZCoobKl9WT+DQFKBvKXovH48rLa+vBnDMR5c
wsJdVdUbY/M7oy7H7mVa1jGSP9ghgTonlmOWmbnnjZwAghLoNB1o83nAdxa5vKNK
EU1CUl7drSMxIpjDcb+Bnz+/o7d3qGpwehEAN03TtqS9CyKqRFo4nes3d0bOChCg
tPAYzOFGJnpqEVxGt7RmDjWP+H++DfazWXreyQQL5f0E4nBE2O9EUpJKxE7sp04a
r+H6O1soWBiws/CLrCQqB632ZG75Cr66AneI8hP8mPZDVPG/xV6IvQL409cpXUki
F0m/LGqUx/xY21/itFAIExXqSVFLJgcUzyfTL9truC4ij3opERf24R4ugNnC66VT
WIecNHr7zytOY4pW0oke7LGZ8t6NKTCj+QZSZEyHahmxso9Rnm5hqy+QyLBJzpl+
JykhbyYT7ecWHXMrwmVp5m6VZfwyTW+ZwszOQGe7mdVTJHZ5BE6+nlQ5N7iIYPs0
0eBuKzWVi97xopwNneGyHJakcldLr5eUspbie6iWGp1Iu0XkxouAwXuBb7a9uDOf
mbIZMY+QY5zBbFMIWmFSg+koMzD5icrU8C6YHLBokmMObwkSSlftoCQn2mjWEZ4/
TMfY1NfQcP3S1nkmWMC5JWPAbTWOBUGvzsHzRdA6cVLElz2xTVkQT8gKSQXv7QGn
tqF1qEtzmjP7XlcHrb4q3liLggbPARztssf8dJE4TwZaAhdzoD2jmfLUx5pTXrHU
xaS04TYG7We/oYtrdNFSTDEiLCN8+U0hVuyjlgtofcnQT8mnq9SRk78FrQ0HICFL
KhNlwLJBPGbQHB06Gl6MuA4AxIZVwuxr7u0mPzYxny3BLHs8Jo4MU9p7N+8+rb/2
brODB59aN1EwsWRer+7cImZqfpg2xIO77Ni5crbyITlB1pY5gm0OwRp6yjKmWTxI
AwYgMUdz1XQ1idG+8ndjGA9tS6kMhG39S6kILQ7tI8VtpuT5b/FR0clllFPcL3hu
Pcx1UDrSoYU0Om0/Qs/BOQJOI62RJx8D+TaijLC8YgiBuc/jydLXK4Lnngcopd8w
JnD2HcRq4EendF8wyruoDz60aNJqYQ+i+KaeRsx/csyARF9ImW/OfWoyIjHSfuW5
28wmu37w4zH7df+2d9MkRxGgKRz5ea+iUbZouJT7JQtRMRVeQqvUVHgOholgRLAo
U2Ui5FaIfrisIJz8M+MiRtpZweAgtWy07P7/FwKyaUVt9XwfJE7JszRZwvW8eyLl
4XZtCLrJLl1l8CYxe4E0tI6+WioBzH+JxjCni9mzkO5sJDinIf8YrCJLtHTyASUC
4GroBwDj1kGxRDMAhXa4JNyVdIUGLt0f2aOjSW6wUPLnBvcl7VdXH8dA8ZzUg3qe
DhxxVWmSjRGQUVqsvEVnxOy3p8dp7QLfXJ29+Ai890hL2qq3VXxeguDrawM4yDdc
6HiGqOVxC3Zgw+aMm6WCtYCBi3v1HFbHU8ZSOVRn7i4UCOWlKsDgH5PIHEFuIsUp
Mrcx4vHSe33GIG7VyuJDea1R+GS062FNyBLtdy6VqJGXW5cvskgYoyGg2j8UMbjX
3wJLVDSz8ykFi46SP2ExD2Wvn7eMgeYbdRnR+/ZySBDXeputZnoRZQB7xtI/rOyZ
rOwo2dGbm8G0tui31c/jq+rmWuQLZl9ztUTvCxXf3mBd/T6qLzIcCHLWHOUqndVT
X88Q1LauhC6ZiBjSmH89sO9a4OO2gtts2LQmu31eSovQsKhlI23e/oj59bKmNpDE
YD0XeIhYBczV3YfSoI9QnvIisI4y5BtnbfHIU6+BYMznWQlTGKqcrCjVTXbMg412
OtF40F7TaazD4MLA0XhWguESDdjf2FOG6DmkVYAiKVXmu4yjEHYhkUGWSEBUn3oZ
ivB6Y+74JoCbWrvJJS9bDNJUO8gRmxPjRsK8gWxAwQUR2s24NjZToNcZwnVICtq6
iG7d0PO30umOeMN7xJ21w1Rfuygc9nR6TP9CiZ6JZMAGRITU8U5MAUQI56/aW6Aj
w3nE5wJ43R6hDdQNDGWIErs4qDM699IUmJspltC2OWXCyTXu8s7dc3nq/m4Wpo//
fzn7NZlzaqzRO9iiV62Y3kP6qqzlxpQDp0aRphJ+YXgiul017pevZCb1vSXeHqmP
q4iHkdenDocbNLo34x4BR0kgOm9JlTXt9o8kYaVZYi9zekX2anQX6/ZhsSca1Xa8
bjsjGM8nAmL6XzpBM7Dwq1Qq34KuerC0YjN/4e7LF3d6+aNcojXiwHZfadE2fpgN
hKL1W94SGD5QTUpdBSvuntOpXe98p3VYzIVf+kgAGeDGuHuvwN+qbyki9JoLyYG2
D9hZY71jSe9qSrnL8Zho1p4w4/fZTLK7tFfs8FrJJfrEDsxmoPJQDOMVpgs+bfRE
oXf8ILGPnq/AfxPCDKW87L8zpNBOeNkJN7oqipdetdjSf4jUd/sSjkXJoL+JEsqb
lYo8Aoh/AWUbfiIzmM4DddmcJgfcq//7Br+D9KGbS3raY3G5ws1yZNRRjSaF8G9G
8weEponyc+Upaj6N6kGGs8vkjhb2C+Zz7qINK4G4hBAmxvltiirpQTtGAt/Q55wP
45TTMtNnpJZC6rNZSEGYMOExWU3roKJ6aOPe5lQXteeLQNtFizuB4d8uPI1wP3vT
QoenVxit3ij+UxrRPjxkIk7g74odUpt9C02/VwaM7l583+2Cp+ptpPTR5LE07lm+
71+gwA1hObP+lCPnefUi+DR858IpwCMmK+vOnubl8nMhqb6dKbFHqLeev6dcu53/
m/iwfz7sJxa+Xl0Gwg4pgV2W45ChwVOXtbY4QmMAx0EEzQn0mSwJyJ2b4h2OvF02
Bmc4aj2yP2CGNiANts7PaLivr0RVtP0NJ/1sSJ0Mx5ZCpsTrw0abZQjhXD2UX1yM
CeXRXodEJOl5lHWQY49HDdnTpS8OUuPncKURMSv4vQD60EeiftOODLYSbuLcZ0LB
3IXHvdxffJAFAibjxwpGygnVBiEAs2f1eq6mX3IX0GR8zpC4vsEqKON3R92obG8N
Yqd98Wclr8xgKHjGGWfs1bT3vqDN4ALMfHuwFks12Y2UT5Pp0jIWLAP/vzd3aaHg
+vlYRyhpxNr6hBB46ZoaX4X63gDbCIP7tYxzOXhAe1qtnjB0wZT7p1IXt6RWHOtM
aCD/AMvOwoTIkju/oPRBgigC8OowaRDZfWcAFwvwQyELsrEENfQvQRehvmi+NeuX
v/BXDBUqyQhTpeigKLaw4UYwcGrr0SD+zfZPr8nJMFG3AxIlPBPPpwdehenE1hnj
LIl02JP3xwSRz8roroSBHyNlTIBzXhHwBnkAZ9D6uiqnfLM+8T1GBf8Y+DlpNMSS
yuBmUq6I/LZ3CNhQCWq1AkdDv4kYjSNMPFk56/zV/Nl5FxPtYYVVrqMla4pJ0w5/
citH6y32onB2yZ5Hejzms+f2BifU+6FjW1CleB4LMGz5FbycpS0qBd2uga4lsCsJ
ThQdztGbgizwZHd9TdNNohoo6AbQ68jN2bxohP79UE7NsjGop4ZM9VJXzHZ9Dlfk
uXsX2lQTBxzOuVqORJvjrZDjmGO3kuG1xZkwUuBfIsSyx6LHYAl+7zk3JIx9t4/v
GtbCGxwg84rWSrgEV9jPkXlPqa6ihzo1ng0XQiB87RPfn4yTyB1atAWe+N8n5kD2
xbwer8IM80SwwT5LNt8rSfq8Twx6r98tckQw1L41NUCQGLGVb15ulCGVjRcqg0eB
v1iYoutzJqXzfwaW0Rwetc4ydo5SE84JFQfAYUSLZWtxIFUfu2mwIwpDR5V0OR9p
VEo3k7EHxsImX1JjSDD39NXC1fW2xmb82mPMRkEx+ZK7X92YjFZ6ARxS4T6ZNrZJ
+vm587vdDKdRnrSCQTS8LNsLV6/NT/bIs6ejr4TgKPBoaVsWj2yOpApVcV2xT1g9
O7XU5DV3rTsuA93r0BvcnrVH/GfOpmgNelWezRaWrMTmaEh8kbyISVBKq6v8KW53
/+wCMpL7kNl+BDEEFH0Q50YaqC2VfVqylVyzWkTYAwkLujTtwgQFbSiGX+y6BcoW
CI1gwyYc1QGITVTP9rXDZknSejncDwuZ7GFTyGZ9wgJCwHBph9wGszBkWA7tBvgR
rCgiNcTQGdQHK9cCGcFQhtx3yN6wFrn7KsZjS2tIQ8NfjAMwsIxm1a9XBE1YLej+
Krt5MiSQHDeoCt7TiFM90D3ti5LswAUNk78QE5fhoZLAky576g0h1EKIH+8bVQPT
95UkHTKXQPnp/vuvXbaaBT7ERmvClcUdu/B8YcVB9/90FCvcdTNl1QpDMz3VhDgy
+0Wnmem1yrnCxm64ZyDZ3bSOfy/E0ZuJsuA6IHziuUec4DFOrgxJmxrR5uuoQXJY
budb9zT2HksCaLPE7f2IqIF3r1RhVdo2WXJZi8DxHhA7Esffd9eUe9+xT2RUq5cw
4OGktfoVRFrST6sINcDH1Ob5OHGx8B0GxVr8w3hK3d9X+tNfkcnLHzYzDetKoEfa
gsv67DE99J6/rL0d57hVWk1BzvYoJd90Sse3922PxufkkIzwh0/wFZJ3/RVAMC+9
C9zJsgHy0xgq+yFDNL1xbloJtF71IKAyafbs/cHrs2eAVQvd2TojfHjReDJBYlhY
+NzGJd55o/+LaJ4ZizZwYZUs3DY1EYPvckSyU0voirGFlBlaL0Ht7+Q7nUNUsyeH
UX6u6LpA9QddAL5NW48ZdoiJ8cFtPOckea0feVb5A8ud+Ms5IcgMwFY1AipmQB+g
WdhR+mdg8uFmxNmOhIbMev4vzdGofH9R8Ehyfu0m+pE70Z3Jlzf3DZR6FTqhcmf8
FgD/ikK3MEBGWr/DrCBC065X9UVU+5/i11Q69aixnc5Uj7w8RoF8L8UpVwZXy0iF
eh+XBc9QD34sy+I1+mIWnVVwLfjr7n29P8wnMeUejrnb8ohbTmW12jndWyUZOYCn
FWLxPYsqiXUB353r/0HTaMKqr/L779Y8wOvyx6Wsx3Q3qis0v0lIM5HQQbyYWd1J
se1wAEHavoNwOmgZews0jkfxcEcLVgm7Sab6+diIrp3d1efjY53gxaeq9C9epBbY
ZlT4IbEmGZAzyxBpDWx7vpePW/+ZlQeck91ok+BOGrYBfa+Fsn3uB2vnsUXZTBLf
YPy3MkZ+A4iW70MwXnIb72p8oRJR/stHzf7smO1NtaQuWdP4FN3tVkcXeeu+haiG
3NmiFRrjBd72swo+6kIRV0waq86mCkwpQsBjA0k54Qr+WlvnTqgoGaDz7AQhvSxS
AyfsEas9dBgRSk7rE8OXZKMnzImYEl0dD0tMZOTFdR6sn81lb3qj2vTfc6aV5gyX
djFUkaoz2cBlXhwjhO5O9bF0G3ShA+kE5zTyePflPxEL59QNqHXP0bjZ4Hc2uOLp
ghfeRDp//BXin8t1DpnjXWUVt+mVPqn70laoT4G6an4fj/nljeNnigShqjkXtCSz
CVhRIIbuNCYHjmZYco65WhP5Y+Xjsa3QtOuRgEugT5upqQTwyNPIZz6a8GfR1eT6
oDBno6o/uKVFsIxQmof3Bbf0KfHQkirDpy9UVCj0ZTf7OAFYiG4xKciDaYW/nRmi
KJuM4Szf+9hTMUvFYIke9REncPHGtzu63rsH2T7ecaiZjVV1f8wC1Lc5ulKUtBW5
IxU7w2Ps52el1qvpeX31cbOUskR8tN/QV8TzYlrQg+MWw4a2v04YL4wXAiZ4PqDN
OcPznDc22cyqLX933QZymfWoKNn8fWsdcZMY5myZFlGmYCrXeRUGyErgrylh/QB8
k5dOblwPsSMjfau6oQtzmf815pjKdX8tF5U91+TUW//TkGfbPeDaGFZJzSiwJQCq
ju53tKbdBC4ccDm4KsphCG/rVOrsgmIkqgfXZqHHIlyavxvpcBgYSsCI44i+bqQr
h0v73FrSXfDMTiE1HoKLXGiKIRuGHG7RKR4g75iAPQyPwUn6cFXbiwFvcTB/S5Bo
ppn7mW2ZXqI+9AMlySkBLe20HJT/QouJiJCCYXHYCxg69oZ/a21/2YlPd/O4ULbp
`pragma protect end_protected
