// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:25:48 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G2sqTLZWXqAtV7hPjdk9B6RRciqmSs6HUZG/IAcSK4WjgAAddiy3Qm+K4UwrQBgM
5xjgJkdil/nos1x7zDiUHjgOLiIs3Y8maNyJqtT9YsjyIygqMgWdDQ5fuPBI4Obx
JCGaHEDCEMrLStez0mbq+K/5foNb84QZGN7bNYaTW3k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 124784)
5m8/PZP8NFqoSqPZSps4fR22Rzp4RlCYoaokNVfTfmUJ6bBBo5cZ10lfQI5u5DS/
Fz9VL0vDUnyLeCMgqgAdK0I2sJx49LD6czkr3rbHx1E0nnQTGvmk7yPAps28F0aI
UxKMdwTvLfsQ7U55B9gHqyu+hCiWzN/8de9ToKds9+uM/dG9qWVyP4aq7wFROmjL
rf8B0uG8lV1c2vuGrW+IPzn2xJoz1PglLIzILrld3mv1hGO4tEUas+ThzegIROGX
ahE9Q0x4EftiD5JP/Xmn6Lc7oJunfRLHU6rkUqXVpOgEFeZU6GvIQJQQKaknnRnv
BELfIiM8YZ9WzFRv5WXXpBKw5OtBAYf9fMMYDm1u8/53M54PIPZhxMhS7CJRxAON
j9PayGqnDEsPPXD4afaNMRtLQD754L1XAunJfUfNI/nxw1vVzyF62OG6ZdG0eSLG
k1wZAhtcDJSCzwKiGMUeAT4pmDoDinzAuQ022mYnjY9GNSW90Ci45km2C4ftMNS/
U21GvD2V6q7xEXQISXKxRdsL8qWaBeWuJM2GL7MGD5CYhEei8Zkf6SqXlaiFnH5+
Zv22LsoPi51sqhombVzjGxymuGncx8ycpBzjIeTn3P6/cRAfXG0EsKlJsS8Icc2m
/IrbRUhG7wxjO+lBn1WEWGwtu7nS1poUebVsng/V+nFE9Aj28AvZ9SElvE2ghNwZ
rAKxBlWfIVcRohuEIre4J596t1Ifu0EcNKnt84xAepV5JCFaWxgV/yawReVbrKFK
e/VosnDirUP0xT4hzP52wSvLQTZYxLsbZGgKdrid6UDXckmODK9Eql1f3wbX+S//
oTSB5w/hc/6P3EOY7RYrDFSytRpIKmywat1qJpmlj2KEMi1uFpuBaM7wnd0Jbp98
FJAC1cMWouL0TSsRPxM8WSDXYXc3Np9SFiqExHMeoZrBD6OvgDObcpENOVl3NZ9R
frvtKrccG8SKqsA4R2Kbc3Fa7BFjZevyshyb2o9uCZBXfo+4zIeb5SeYeQO0UtqI
MRFyveT6Xng2GrE/xms4kcNPEOQlh7oaUQ8D2fo0QHkRycocGbdpQEt47Kw0Gsl5
2Un1VGCnEE6ikmhMFrz2FGlJ3k4zswC7hJkQ2XiTra2G+jN4EMWvfdb3vzYnFImY
/31KJ67PfRci4vWVD205Wob3lMs0tnOQnaZDYRU6RrADQiqFs1Uh0b8kL48wdTIz
VPUOns/tQvyMimx4gegDy9nUVtZ7EsUd8o1fCTUHLU6Uo4j8Xw8sWNIcvVqwzqp6
yeBPGkKlhbs7TKCa9Wm26k7scUEJ4P7ZzPBTv24tfns7clTmJ54m3/aZbgjHMNX5
VrqJJDem0c6M19jzFTV1HIEPdWPi6DkVvGe3rxrQhBHbGBk2BpJJOv0ysnVCNDNQ
K+vuvpmbQnvZYVBKdJ6l5nmt26Z6zMflP2ZIB3wJL8xvZyP96oe7fgpFW/lvaz55
8pByV+ubeh0PRe540Ne8b72QCN5MJVHynQfHjw8JJQrRDzFp5UOzNeFNQWtpaJ20
Y81YCD0FKE1iAloKYB1wMKaPiaphnE4sweXGvM++YEGiDbjz0UbGxAuOdKdqhzNU
0uz4whXm4kHZ/hKsK8fQBndNetDpWX/pi3iLh//YLF4o7+hSSoKDRI0mDHfMXPxT
C4QaQ2cVp6dkVkyw8Zut5MGryawKx2mrGGPiX9mN6y6ahZ90kOzHaFHr4nuyHHFN
TrNZfrcHWXnsn79DgVDzl7MsfF7/wZZu3td7blGhGOoWTw5kzwQ0LZi1Cn58kYzn
SgkbrR8iJ2J77NQ9kFlV8JDuhPbDeJDVUhSo3jI33RJ2C9ajijk2G/5HS2idMZ6p
ZMhivVKNahTI27fYELnnHwC9fp90Y1RpHpjq0jQ2iKIFDrjSN4JNmYjq5XSZHw5b
VMRuTvJSbElyI0VinkRaoPBlbgjmTOpQTNpArkFhyDmBe28dPbqATJCMRxLKDA0B
HvWxi7UnIBRR8MTAYUrIjDD9/Fh6vokze+kOJPfPXKMn1kXptbuvDunyy4Rqh+v6
eresB1C4YgK+sYauwHTJSttu9uDkSp65sCPu/EbSHIZ3nopekS0dJ76upk8cU2DY
e4sS2ocb2Y9efd3DRKIyjd4/Mr5wa+UFwkwj2A6BOS26MiJdV501Flwuqo568Xa7
3ZDkf5lxY3yGFXoK5l2zYWSxYuT7B8E6HPd+MjAkjX6qfcqQr/qVE+GanCWK2Wuu
1hOjVAMsIklCMMH3P5q6TgFaiBBpTqjq8PJPlwNSk2AnFHRLob7/B0hUXY6iI17v
Rb9ZslMKQmwga+OFUwWWHsarCpG2TEsP1KJlaJrtvwpSd7FXfzOxe66O2vkuu200
pkDRwUNxTI0uMZQdybXRq2B2CG9+GbadtacnUGDtqX2dOkwFrRkgctFzqWtCGzrI
cT6201BLXuH2UfvwjPaCIEqmG2iCYol6dmOojOSt0pBcpeNDimHDd7JL4pIcqYDU
yAQBlq4W/pAIKqrxOVs1sFZk6+w/9LtpYqDqjZXjztSsFibT7zNuNR3fgrAbXiPl
D9ULSUk19jVU7bJSjU+xBFOOvobuvLTNDKQNaQ8F6l90FWuPZZK6mQaAxHtYb/Nv
j1XdlbK2swY0JGF+sTdO5LaNvOdGOWSymlK/Ww7Y6m7V04WVPGpDWrGvUY9sYxoa
LFc83sjoY6NyW9X0Zvjl02cqEL9olGajJOQLUX7FppHV+UNpuYqQaGNlsEggON4T
4mFlrwxLdxqyyPZZxgtqgDB5r3oYqDMzwQmil8oJLRirw6wf8H4UFyZcSsqHRj92
OVwZnVssIxHMFQEofdV7j3Gf8PkmRkwpmduUDRmILJyO6x+X7wMYjB4a3gPMhvhs
phfFzdC9zdVEzLUewTdEMtZy6J+d/22H03bZY8lrjTm9MDdQGg46GyfZdRkQHCeh
33/KCuXnfi70lWOcY9kdRH1ahDW+fYnq7u8/PyEpJUOB6uyQ9EzF+lBIxQaoiS7j
cOwDNbipJqWcNHpJvJutaIcULBCTJdCZNQmLsrZJ7zs5FnCLD4IOjsl0ce7wc5KK
qIDP3Jg5UtuxPWUcknUUpVgqgrFIJekBnDDc9fLFdUd2s85oeUKsA9XrS/ouSamf
iBy1YcVPZmKmfR/RsHBUPMNn+YazkecPfrZC4xdPyIHOYByZ7e8t081Xh2lQTDex
mlPoUCflBbctGOn5Eag6ulAXF06G1s4AO0EptDaDRBnkFRfGyuh5Ifo4D50iFlBb
r4MZWjLFR2bp9of4zxNVzXl3bSDcqOg/YrdcRwp+Ko1x/xSvL3srOVvoWteS7DIj
w+khFdseP3fVRFef9zDcAfNhGYVyog2ciI/iEZxe8ntBxIjd6q6KtTmAr64Bk3yd
HnJyeebcNtfSI6L90t4k8yT0CoB6jYcJhLvqXPKZI7HQBOjdGoNAtYgIyl86fDJM
ntLci7OPT8Kk2bd83Jlej6oDSIfjxGk6zTB++Jwyul86f6quEqojUOIYmKXuK3+t
ZchYSRNUeh3zZuTb/bn2q6AxODnO2kp5b2JCMssZzPXwYzAv8xyTaPDF8pyce7hL
SxP1WSchutBMDCzdDUGpLvFP/7jjOXoaMe6MJ7JaEVLAtaKGVsxpFMxAbwdRYM+x
LoBc1wdsq2Dk+1w2zkOM4kZoEwlttCmieAJzM5VBolxq0MzKIbOoQEtxxLfNOZ2c
79LEpF22bLUOlJM1y/cGrbGMdSKVcY1P2NNrXEI8su4yy/EW1oYmcttnzB6jrtly
i+9Zj3jKQSVfLq/oKJHFDDkU0Msw9g9iuVOclY3yrh7b4RmcWc+VHD1IEPSCkSTR
W7bx26FuMabnT629k4GWXwhNqbFxVKbRbb6MuciucQUnbcLrmpPeKQU7ygWZzgbX
S6JufrwzCp88tkCnEm1hnOOyiBcmGD3coBLyZxB8VOwJ5XJPtxn6TUU8jAQidWlV
pXcraIH1J4jApyHHpGlSVJdEFYI53/PBhM2GQkvhjQyBbwOTfJN+Hf4sfatxUqe9
j9WyeC/wz6ICoexnVVxNbcVRoCQ60SwX6SWt+bGFqTal4yz9LboFHyyraw7xJIOx
xE05Xl/qrkpAUQOlthKToyaTtCKmytirYA3ALx6ispviFWZzqTEv0qvoLJuVxhDb
ryl8WFJW4ELlypkg+iMDAO1JdWJ6P3G2+0xHI7O+3T+1rw+qjawwIz3WhGKPfK/y
UJNZU3kRlyz0V2kJtw2MOOcwam1HyyAw8HKw2f70ME4kWw62D4b9RMJzZOJ33FtX
gOFgrENsCfGqlrNA9gf/5pxfgGtwCTOBhwJdenuUNA7z8jvSZGRIG4LaNjaTDiQr
+ScMzBE+c/782+qC6X7a/37+5qHOh2vFwi8q3NfR0uUlm+sMyKHlryzCbWu/nS1j
+i1a8Vi3YOKgdWeRb7lGtSMPHyBymPruqNhxuhTZHAynBQH6G8qyeK8wq8DdNMWd
wl9SFnzhiBnmowUEoemTdOENHWUIk4jXI6/mQzVLNLwWQm+gNgZbWJimXZmXUf+x
WrFo6c24ug/6E3WJXcfRhQL8aDFOa2AuXYJkHhedxolEv88z/lSwc+BvqzxmhBGS
gv3kwWQX5B8kCxOZ0cldjKZq6AZMFwRTO7E51v4/YVCL455zaGvL0s81ALC7o9wO
qPSW7B7Ot6TTBLO+ysVOugCmV7LBA7js0UnTzKuUFsYd+9wjmyZMjAYxCHDJuhfe
H4Inbto1FlOxJPf098heFtErpO08n694AIkWerlu5ZG6SRW+1jQLwBe/ak04MbCU
TqgEfOeSsQs47MbATruLss4sg4QlUXMRAPG1m+wngelQAZtTCFPbgiRYng6y/Rbj
/ELwq5yEut5UBq0A3qAEhKio7fxjJRnbe1Ujvqlcq5wsP0A4GNPlGO4Ub7DhP8Ig
cbZgFOz7JY3zRV3HZ3UPwB3Zc5vFaf0JqLJhM64xe4gDv3vXuWKKgoG0tGpxSsWG
OD3+YCNkzxjFqifEbWUNXUhA2mgAxbtwJ4IUXOuV8TCxO7P7nmVQ+k5IM0YzcvOC
e2cKywEQV6SaSDK7/7cAoBGLwoVDN05pxlSXfkPXUY5bZrd6T7jGidOuWMIOp7sQ
DfKzVYpFAuf+sTdqt6Y6KkxqY37QqgVdOi+p6mcANFEKSXNgGOtdgbVQ6dMs5Y7y
ifqLDvk35uvTtvqRHBnCTAlj98h+WU8UnLnps/9PMIfqyZV8Xi7ED0msOQOiHKRT
4Wspylaj1f513d+9xeY4PxKPGsrRsY8arQ0w4I1PC1hATRLP9T8Wg7/jmDt+XEZ4
5jXgsaQVMLrJcML0FhTMUa2iPCH4HRKapg493BcQfQhy+6KnH/vWmqzSNydNBs4Y
8Z3P4lgxUKK6+u46VpGu6S8NabBUQRYidCBCZBZN+WSD38z/9z9++gtCex/PsDIS
QKWKP5fnlCgKN7PVlM4h2yL0S/q8YLJluXckNYez4Xv0k2eJIkXJLf0PIfpSKLSW
c8llHtz/k6pNgeTVf5nJtSyu4Nc4pUiBVyOnwqIMBBj7zNvMvM1MQ7vWmbvzC9Ht
FpJxuWgyvCNiOCVlgubNAvktqKv0mZBFECZJmjJNkguHqDGCipEWRvWvciUTpmgn
fKPaaqik06I4AACuynmCwapJvsalgfd2sVreQcwOkXVq70NQoBUj+Fp9TTRzdDee
zQyL5eoUGBCezzV9W/ilCX43PZTolLSXjLyT518YgKlAcrD3ZStYyhvV3lRZ5XWs
2lQC3oLLppS3r6M9vz1y8eBJbYuCO8A/QhbWkriSsQxYaaN74+zJ6mddW1zBr6CU
0UGfZiorsdSs9D5QqhF498WbPXY8qNm90jSdPfIks3sSZp5tCwt0cE8Zll/LAeD8
25yV9LMoN85FCVDJDHZcERGfjotVe+LHOEPZ4u0/26gR521NVCIn/gxdnYu1VfDv
D+efyyhlhS1qXRoF9NZrruTPVtKyWFoic76gfaG2d4Uomo1fdFENPxr5rR2tH0K5
dwL8UxTubC5bkICvblswmtDq3K9kCUyIpP2INFOaz4aLDCjL3JGMZGxpFxc/Swo0
zFG7b49jDiiEgfWtukQGIART+QiDu/9RX74ukZi7fuFy115VeaxiEs+Vt/ZKmGFQ
S/RjykYKR3yhH/REJLiEO6hzo5WZaFf2fnqLBDOm1z69q1FlENNTxc2UH3s6aoql
LODbOPzNa0lJjy71Wj8wkjtVE4yGeXE7MvVjyf8Ds2oqhzR8AbzzT89flndy8Uab
dyg1T4RODcd7TfEAaIdSrjjLTgxAqqFomi11RruaJUxMCYuAZ4gNC+48Pu7ZwD6j
y9FYURkeamaco8N1XGmjVZbGvz1q4NonKBUg10f7bv5ivGZqvLHreNBlMExSt//Y
2CPrq2siwlP8uO0xNvyKekXmbaVJSI8R1drNWz0uLBo4u21zoNEj3xl8ctseLjyl
h5pnSJDU2bzg6gprjXXWax6sZ/+BhBfQNBkLPgHjdD9gN3mFdordwPfhivrqVW8K
XvDaV0ttvLcV2eSLkKBisVrBMxFcP40wdX1OknSXvCTLIroNtDTdYBta5esyuQi0
6MHRmzxv+OwoAk7Gyl50WzrmyHcuPr2cBxZdcvIJKqCd55uSESBG1xNaYdAU5OUi
qJUmt/nILmCRJbuyKnae230ncNiSycaDnglvULNAFl4KWP1T38P9DI1t6Grbh6Xm
JmIzVA4ErcEXWVjXN9r8JYHl6R4PCLw7Wd8b/MPnFmYAqixeezZFZATNGpPTanLU
Y/LAugfaHmcCKVq3MQwe6g0F3aCRnwc/RfM5YrkVALxXgLJUd/p7q0bGh92iTs5C
09fWLJWMw+UH2T3PJxrM3k/owLIQTOFigK38lq8eI53c8i5GhKBdCAXkvIDSmx0N
M3qrKcgKo6Wbh8/HVcnxlekU/XRmhi1niB+Gq1mHPr0iKfzRv/Hg7/jeiJ8UVz0l
qxk0KQSlqiZIbnKWq2efmeSjB89cG6juN/YRcn+EJd5iAhClSgv4uv9+hSnzAFwG
W44rOMePRwbBvM6UNRdkD93AN2eypbQdH70DFlOr7IJLL+WipGCTdt9XoWIKv4eN
LDf6PR9JEC5mT5B8hKZYuVaOc/oE8aers6sWRCq58h3LqF6HkZ4Xg/P9myF8F0NT
zwWInIGO5CcaHfGdZGKceEBdq30lgTtj3PcedeQ3dgAc+ZmpTTiUhl4SY0YPDnoC
BsrsS1kNjcqGxSmdOABZDeUT44cU6YyzUqyIowyKCp9EfGmctShG0FbLYsYue14J
XhVRrjmZhnb9BLki4Y11xtLqmV4GkmCtIEMwVpjLPuzHN/Jtz60na7QDLCNPJ991
R8SYOE3/Pn6oha+fJahPfFa2KnojhV+6MWk2TazfQEevp78FrQ+MUNZV9xalIq38
o0KBIrY1wo6UlfLdjJwYbqPLadhUT1uf8+73R6EhAOECJQwHcc4o0oTqCuX8kqDW
BH0cFqJstGWhsw4KRlixe0wZIleTgRwuah8yCENV0MXfkmoZ2uk3ARUtpdsJsRba
rw4Gy76kYORETYmTMirRidGHg5qb+HROE/DPTNqlZ0+sc7hOv3farNAaWRq6Ieqq
EEmKhdtLQ4gbdkvcuN/lepe1dEDRAufxGuAB/aYzOB04F+I3dzpyiSet4bS5NOta
waj4Aq0ckSGRhnlDhU9kCorxmasqtyEsJwvuMzaoqprJZvXeeQHItVWjPFirByJI
cDvxGZu8PJZlfDPzdl1KudOmDgaXDFVd3+paGctQkgpnR74+CA5q6V8iVBCw81VI
ZpKo+ZaJO5WOxlmbmg98BD6GZaGGGR0hEA9MjYFzYsBBDT3b9cLsx3JnUUn6+kRB
9WFRP34EbWmIdHkhFux+P19nCLuheW3WcbW01XsZ7PFNk9E6T7UdYJ12FlA95ZWq
0bUCUUXyWSybb44PD90PDsb9AmIjHZtM4ytliYzyXsz6ZxGNegCPh3TEfxiGtNft
sbcaIx9HjVVoefEAFuaIl/PyehZp5WXnN8Vdq1+v1cWZ+TjRUSK3/DSbFcPMTrk5
3L2raREL1eA8lWnrwehyh3LiyF3OrPpzadU+vshbI1mc+Y9oxTD4G/0blUDmCP16
Hn6kUBqHHFGPvoS+OHDDJGx9wS7H9Hf72E6NkUC+tUSMDPtUAlrXdtXmaHbP4Hh4
CeF2f0ajCxhah49NaTBeo1POvO8XST0PKdWq65TStpErgtNVrvoCDXpaonQy45mx
BMuYt1BoQnX/5Fj+wykTN3UZJONVAYbY5lHe8BftiCflCaukFvkJ3kjF2SllCEap
eAbORqHPPk5i7BdFqBZruVv1sa+9aa1+gKQukQitPl8E+oUKHbdXX3E+cCS8VhIM
1DNM7jZyBrBJ6ipZJowdepvZc82hEY4g4ChvglwMHh8EkI6lhxcBozU+1cYdOMNa
pPVuC3gzn1wOSjz208r+bfuY5yP+kyj6LzVuhBDWH0A0jQJ4+LUp2uqQJZjSJ7v6
uS+y3qGiNn43kZsE2en2oAQKbg6bVGSvPLuAvTvogiM0YOu2PaGB4cDtXdFammwC
VNBpsu+edA4xd7BMXpxmEElHRW71vJGwDjmIPrWde2RiCpt66cBXyYEGsHrbgo2n
0GKHHdMahnn75ue6Va1kt8JFPaWGgghDL006VK4LvOvj9jvAe+kHVX77xNkCW55G
PkpWseydUxOZEr5lRrdi7m6CyQRTfG8QBaXJXr8mO9Ed2ZgeWVlgZT/cduabHWXT
rf43EUwHVDQZz5F8l97HdvmlzCAZcWJsmKNucsFqWpT1t2AVSMCKj9XmINWdaSKT
Z5ffYbppkdS4wNM+WduIGE7BI6Fs+wmYsfWFS7G7mbvuXcA8uy0Z1PXZf7CvJHWr
yrHZC9zdmA0opMtfqvZOTQANgKvPXR9IB0DUZ0yYe9bat0s0UPpUKDYox3qze0pU
Jpjw48teNjxGLr+JYdRVrKIMBMdvTq7NmrX8maVzMvveouy8GBdvKS+aATgg1B/q
mZefWJHFzssPSELzJ/YKr4AUOO5hO9a2eu+PNQgWYnzFIBXnGxkfJzElvP7PjCls
NYhXZk4u1YGWxyvyv2sghyMHRRRc9Q5ZQ31vTUVA+/BIYZe3dj8BWYWGxWXr03Av
H9CmhlZHDt9ETm1vfzlgaQsEvjfdhMboFxy5POSKbpxz9uPDlNQ1lRgjXDqLnkcX
uF+aTll1QWVYJKu7f219rSSKV/8yhgqccnvlc/UkFfcJr7GMQiMj7jIMH5XhpTwS
zzIpytgs1tm+XP+hH1elVdvlUNFx4bWkUUjrfR4gk+PRdpmFZ41TJM/UhgGofgAt
LJMeZ+CBliaYaHiyHhGwVFxxFgtiqjgVpaS28t+epfQH/thKD+ltPqOykotwosqb
ylCkGw7QcMhh6KvbDO4wZiAyhL1bwHegFA0xluFJAnCIGMcVsdQjI3FPZnybWaV+
GXq2dCG5vrLAyT8GgKC1WyH+n1qsRprXu5ufAQ5n8C7sIkzRLlL5hHB9lXH6A2MD
hYYoIUVaEkLuqQNBVLrcbWswAUJ3re0Hi70FMq+CI4uZvRiFA3tQC6pBZiw5D+uX
IPXo+6INBxRDEY8RKlZtB81y3YXOG/gwPtYieaTY+RT7fU+Tu8XicsgGPKxtddpf
EbodqCmLRjyh0kSw5Ay+Kw8wNbMns983MiIKEu2MmpSoG4g+A5zGD8Gx+7+mjXtS
PbTs+/woml8EXNE+9JjEIVFogEcvgF0mRIRr53nEa5CJ2ZlA+q59A3Q6Wyh45lJw
EhNqjLDaqkXUa55FGSGqI1u3/QOvF+ro2L7bXlIDxoQZdiTVuvOO1tAaenDeSXEe
/VhnKHYjCinhppgp5JqRljlNyEbUKxLX3+PVkBIsBGFT5LntCp6VPqp1NOvDLZxV
Kf24TRywViGSp/ARTYnvzRZmCAwMVOf2joF8yWqq4s2Dg3AawJ4bPiHMCfr9tybu
jyssa/pq19e4TeGflV9Zw0qyhnRL+Cj6Uq/4x6yqc3jIh75nj6EllGtp3vEL1NRg
OyuOqPOWBAEFAPfdM8nmRGhDQ4p3ftBfbZAPbwRzdYF83sz+mKYB/2sMXvqZKqYS
k0Jj0cKN42eimmFJk2txX3yHYs2oGLeyqi4yzjzG+yPkYsmH48P+lUrKmqJ+B3so
6wu7/zUC/ROdgpB/RB/rjc6mbdwMzOImQp/4OgNFK3t7YLUD1D6iDhK9GsWjHyQI
nafnkoXiUGvOYZaANMVHIZFlwyRNgzgXx1br0l0vItDzztcK89JAHbzJFd6st2vI
v9GzD9vnl42Nkovyr8ltFo0xwgWwXNOLK/UvGUedN4F+1kwHe0Zd4kwPrMxZ2amb
RvT9KhlNjiDG0dmrReW+1XeQiExuw+pAtij2ocnzArVKih5/CWjeUlDGkYE4pZ/4
7nu766Q9R0rOGQzrNXbM+gv5pzKaWNNyMTYrIs+qngCOlRP8N8LQN89sxFWQ9oRE
PdhL/M+Je31mwfmiWn0VIK9BzFZu15gGD8EZJr6i6DghD4vtNHXyYf3lVFdg31MZ
1lyELXt3vOHBGwXVi++C5NCTE9Gr+lFYul8EO8PFBvEF3qwgb/XCadRUBTKV/j0v
g7jXQ6KVdXr1Dxakz18dJRCMh6SY6sEQDOSYsF+HP2eVzS8EkGOz1h3D7EjTkBMd
/cGxQi4yXt73XR4ouQ6+qWKzL96Db+5EjrBUp4Gj7eoWhCcNTwhmIsQUdDqL/hVM
hfd4SNbeguWxAG704kCqlmx0eyghjSBZDYoT0Z9mbER7ZZYQd0T2N76PhScH1IQi
WC/jLjA0nDvSvoaHCKjZmrDfyLU/rWqQb1qdqB6XJaNLtflxI/Cv//U8C+90PzeM
LM2RmIcxNZ6K/5trqUeiqFOfttlRquqvC6Y9INjoZwaNSm1VQnMttT5gphY/YUiP
HFjX155P6eUYIbQwELquBbFegDiXm6/3JjMq9qvxFuw14WvYmDaTMaj4G0RnJc3S
H68dMmiWhenga2hbgsbU/RNBICJMfbNjdQZf3cvBEiaPab15hAWI5gqjavMUpV9x
8jyp29pOXQ9wmr6VdHwTsEzHL0fw+BTMWaLcjbQY22hTSAAe3+pCY3de6r03t5wZ
RE8S73mBU8q24zzidCuORRZEHDt/NnYoUXE5fZcV+ktsC+m/Sv9cbMDt9tyMhlLf
QMqQYcndTJNlqQ++xDRibHjTE8Zo9h/qI6PtiRRN5scKTpIQoHPm9925TXPey4FD
mS15UaC7Kl/z9CiOz7OUtUExwAygc/AUNKoMH4lvyfM5gL8KIHTRMZk2sd6gp0WU
TZmfvx3QlyRbfWe1jtKRds1mdC6U1gupsOvYfElsIyDiMtCECDSrzd5FTiN/jUq3
2FgBCrl4yr8JwnqV5o21Gs1ozKGXmpRoc1g9UNeFoe8+a4SGFZTSn4pA8KANHwar
byYa04N+BEyBFHsD98zZ1Mv3pY6ydQDurk1Nex2un49I8c5HCk0YmaO9tYmLAsye
Dt75PxhVYNvpL6CQo0dfI+WhlIHDmP1no9BEaVWfig/2bzlVW4h9B1J9uGihaQ9l
BBSSxfO5VCRogtRAVinjjn/YHBox80PcsOL4Rzkek8Vtvq2I2MtAECm2Anf2o8cR
grpH5oAl/GB4vIPszbIIoyt2uZVFeCyzu5AudPnNb8hx5Qq+oSuNTQuDnc1yIsPj
yIfrpJWvDszwQhYT7ne2IqBSph4YW77+qEMjlODzTTyynQ+mi1cVM4g7L+uoBxKy
tQf/uyUajUdlLdMbtfH1LDT595R88+ynxETJvR0/50NU31Nnj0VtGCww1W2WEzMp
xzM9G5Q8DLLXNnfsrn9MmE7Ms2gwJtul4S5ekpSVd/oB7c6uaysDTQcD8G/QKZ/X
tnkj398o0CuE+92GKRQQ1mJtO+chHPc2pH/tPIL/e/SpveupXn9a4TTJVAYmXecW
ZceAfQVBE0weTkTGlLJaWMmIK4y4fcBc0zJU/3n9hUw/eqwe1pX7nfTfiprHEcqz
9z07qAK3wSJkj/ETJsPeK0/3Z+/Tfin/4fSze5ut/ulEMpu2eAOr2pZcdxdTRHK3
XmKJNMu/xCo6IPEbuK0mtSFj16vbmUjKzQizVhI0/qZkHj09yPjr8cmINxjVNtix
y4ltS+BWZBuf6cyoeOSywPM9NAw2Epn0gtPuNGlsd/c8TqzC/NBxVhh5uok+CM3E
rKNOADU1tgJhPfZbzem8CNQDgxvItBIKtYcU8+2sa4qj5YBMYrSJ0zy8XZFl/9KM
0Myey10o0GyG+1xJZtws//RJch/RF5IzqyYKz6q0PTizQxhfs6mL6ubafUIrO7xf
vrtIS+LvKpVJXVei0NMol8pQSLc+93bkh6+4pAegXapONogculh2f5ttjN4Kj9oA
umRxTEOL3po5Or2sCIhI+YnTRasTCZZeC4G1oP6Euo4vheZzhiMy4V0XIFvMEcj3
kP2/UvsmMSeFEh5yK/SWRmTzr1WsuFXmLKD9lS0qk+ZvamNh4ZdsYIpsRdKkHEF+
sgMMVVMIHDkqr9zaLXbVRHfW1dL8aCclZ+Ma6Bd6d7zwYgRY9P6KxUiFCWlM1o3j
6mGqBURgQtFr7gkUwyKugIoWNZDkrFTx0DkHCuM+oilYiaMjtPIIE61Jj7cBPvaX
lIURJQ+93lEkel7bIhJdfImGznBL/A57Dfh/Cmcjv+fr0PcjpFUFjHfRkbpDIJHG
5FB/zhcw4qEh22mwYrk9acP1tqH+6CjAJOUG9JbcaGe2LNwwrrmCRCr+dbo68qkA
8xW2bzN9MfxRCo1TZL7llGOrK4cIndkZuuiSiOPeVF8tN4h3VtGOCXJ89bHbh8mJ
FpKE1xyzSMsfIcNlmoW77qp/H2O/4bbm8QWE1TM58fW0tEm4GQ+2cj3CkssZUuNh
0ctBUGRmkWOXjezqmzCtujnNi9h+JHuot7bJerb0tY4zRsTuWCrMg9tPamyfPmNn
25XI0RM9TG/0sJVHIBiTvWwMJrtegCtqhlzZif8en8Fttlk0FZZWyNx5wcY3ds49
syBZzZtUm9CEDlQ5aSc4uG0brtdgKexs/cZWIQGjMsYdktlan7R3xNj6FaBYSX3u
eAC3l8TVVsdQRWR4Xe+VXf5LBl30ZTbOXYZE9V0cXkqlQmx7LJfJJDGg+bYBrNkS
lACPwxZzV6dYUZk3G9ahqOkRbYy0M76Fx7L6ddSZTpivPTcgXaHnIKak1aSKFS4x
W/u5fNNVY3R+0EKieAYlWIVaU7hJvAuFss1yAf2EzOTTZJ0e8ic6N0CJWgMh8Eoa
MD3oFAyQFu2KR0YMmWlFm461o+wowStpaGV6b1/vpX6Gd3Sd/Tx9XsWCvd37Ejf6
NdJZZCNw5KYtP8bu0kceChO13LlEB6oOqmt2sCvStrRIjfiy1AfJNFc89pEUbba5
kv1EVa9Pv9LOjOikxkxArB50hMeIxZt00AQlplBcUaMb0G4ziN5j9SZCy0v6QIAC
wjyFbWxBN2gZapbP0dJn+FxMFSKbPVb9aXqIAJE+BDr5yyONyvAR4rDyvi3rvNXb
cedF6VM4EJ9d8MadcebMezxA09jPYSFig8P1dWICCT6daQ18j0JdbbqdlKFEhQWT
L2eWvNT95iWIVLW7NoabwK10IV2ZPIuZvFO32TaZ4EKiSE1c0jscWvJC/IRRzbCb
FNiIW8YVn0oM6/+eznR9XXTze26bj4EXc5zmAreh4PJoUdnEc/EB/2bw1HHJKWwo
SWK3WIns3IcVoQ2K0/T4sxOzs1l/K923clJEeHL0esQttG+5XGtE/Ez1NgnfBpPJ
RrdC0m7Rgzri1zTGtx7J4QV9og/iRrBNrGGf5Ls6F9uESD+tmEIimDn3zJPc4pHK
4it+rUskQ5s7WT5nL88ekUxJpZ28FxR5EzQvrJ7rSG0yW3Jx6fizsyMd7dFTyAOB
rnxnQFV8ZAZYrJWLyerSHYuEnigDbdoqcWANBBu7H62rK4d2BEpAru8er3bS1WaD
RO/JPlGhWGmSWfOvNKbDLWd3B//G6yHjtBiPykKryuRmnnGBkoXbeUpZ7VznqVGP
+Eb85Rsv74nnwg0ZZp4gb9MPZZyqPAZk4F+0K9L6TLRN+llEyX2r+CjH+6tYHZqX
A872HCesFwiBve2DcOBbk6zTsU4PcOItqBZymRdBacTLY9TwBIsgL4FdhY06X0X9
kL8ZB8TLiLZjx+9GjHXvVvysnYqCanH3sOwaehGfjsCv8qV6KxjpnJB5qaQ80ysA
gyJywuSosHAD14xOFpdxWZPiihFd4n2FqDmVOBPXsnxQ5ITS8Z74Fq0JA+LLbTlQ
GWV48i2zA3GDA/Zb4X+eygTKnGvXcT2U2kGMGmpVL6RDBoOZ4nCSSzecC3KrdEdj
w9SNLvnpDjtAXwozeiWqFTz3nJf+4+nsrJUgZpz3r+MSBiZv5D3hA1Jc4871pQBh
OoNAdw0Utr3XvdHb5IAJbUOQe4lvyFsV7uLTcdqIp2r5A66xr3ROwvVHB3Hn58zG
aUIZxKaODsTt2EXs86sl9yX88FWEOJmJCsW7uRZ/TcB9cx9bT5HQQrNze3z3/0nq
vp0wv1zTiGagB+b1Um0PiuPDx3rcFxUfhoeqabZFd40Yf46b1QxrZvvkn9SUyNLB
QbiB0p9ymIynx5FU2wTzavGQ4qyV+SmzE1rUoQEs69oKgResIjjLRbFlpY+RLVzw
120DwMl8ANdFM+yg8eDrt7pkpwu/u/46/3P1Cw0+91jBDQ1/mTWzBnWPn5R/PNIk
7sIb4E/4kPtqIAdmBr2ArjKBUj+QV4d1IV/YNX1RbGm2StD6JwPtbflquJu1mDFn
+V4/0IXAZ7sCU9Xd5A98cq2RfbdhUjuSqARw5dV6JIbHhKEdaUWa3N8HdJzoIqE+
8GJYaLbCZGszLG/NvjcBWAe0X17utyGZTwjKk2912w56ObE2Cj1Us8jS8HNCThGg
8PKe3wR/Vas49uJ+lMSGKqd9NkSvvjYSH3l8677wjBytTKGWLu5od1Uogqrp1nOs
S+K9PvkyL4+JKf23/N4Ku1UOGN6K4/dQBETphGBpQ7njLMVLaV/Ihl8gXNKSkT4b
VyIwL7neMgbGdzOwOcLJy/bJ7TJ7uWChRN2iMJLaFzMxcx8IclgD4WKXFg5/dvnE
CU7BINVy7DaspCo96S3QsDAYn8S+O7hiu9+6s10Fxv7O2nGsQkaLBvaPMiExMW33
qmP8oqNkAcD/bbnhBkr5TzDCoov7F4fRjGDIpoCWu4TmmQJZxFoFD/Zjw3o2Eb7H
FlZ0W4DzAOr5MCKFCTEx5jeuDWYjx6b3AE2AWo5H23ebNikfoszKaumESg72FQca
NP9ZIG6cMd5h1w0x14TwSEU5YtFyXjRMRzMoAKXUd1vgdN5w7q66tBCDLsP5H4Z2
aq598l+zGrk1DYLRKFELCvheYdL5+Jp04bbu83gq72RLcrE+4pmcdfGCcKRr8K0B
DHGgzAwHKZCpgCrZF9uT3Y7ZTq53Lp54SvCNDa8ZIv5Pl5M/HGszZRuPco0kzlRQ
c4X8P17/ZW4gDD35EluFY6FrgCF1qAGoPqcCw+COQDaGWO1RWfTmOWggtWjwqZaU
Noot5AjXQpIKw+tYuc0c85tpa16odYcRbejwzMtadjZVPwYMp1lopSrvzB5gqcok
s0ajPkfp0yjL7q60hcz0eNtsyBIW5Lt6pKUmGKafXtImSEwacrhjahtkd4pYWq/D
gd9NDrw/rHXZkMxsuaIn6teJUz2DJWolZkcsfu7Jb9VzZnODfF1xeGs5hmP5W1F1
xpS6bfd8aSV1NNS0Pp1sp4e3jXtFjHNNK1Ng4ZNfOBE+fDbxICS2x/GA+jCmrDub
IjJwgUI8tsGu3GHSmMBvV7XW6+NPKhe1Vhknx1ouk+DcXQS6BkdiYrwK7o15HG3d
b543LeAVCx772Glfxdobjrkvw1gBsEZ0T952JC19AasWRqTFtvPz1ZJYKSZtQM4N
fwW9jFJTj2Sv5veb4hDmwdVCSKRCmBj/aUIRSE667R2nPwXe7QUCpig6Q/OzXOwx
Ds6KCHIxs/VdhQxXfHcHSEh+CpgLDkQ6kkyRIkpEJ63ozNe/Ju5u0Y37btS2xN7u
wnSx2kZFpycuzKCzqFFED7PTdUq1/3XY/DORWChbtdS5j6bKLoFxTqhRGXPbtjqy
PDJfm16qU2Zj+nzrRLgOi6EAUm4z7dxZMBsiwAJKEHyBhDUxQeBissU4FNmG9l3j
19wZC9DS0Fv2Es9HgCyNq5rh3gCHZn8uKfXuYVnP6G00rKT7z6PIb5nuuqb1OaQY
rtr60PKzr3RLDJKTupQv2LByrqPO0IIWobPVOBO1H88ue/biWatofcNWM0elEtrR
zOTrcbAAoRSn0zxrwGBXc5+hyCnSSrElTQMXWBwZjRxPoRMwwgj+Ov2H0hFz0vHa
Rkgs4XXiql9ra8QS3Whl5xwRvKUxgefjoFYOse/E63VJE0+HyezqP8V95wO8lbB9
OqW+6EdD89sW5pik12w7KaqKW435rXTGIFFDLlR9JHkQub2oELNKX3ECYuD2hHic
uvAUPvhJW8XlssRpjef0ePKsFE9yudd6h7xhiHDYmOCH/JrrREl0UPur7tWVeHFC
wIz6gCVbzWlPDDKGqvVjXMMuWPQRuzrpqHqb3DtVH7EIeHIl+aesOM8Sb3t++35/
6OCNvb3TyXH+UZKd3XmYXuLJB6SEoGaQYErD7JA8q6V9o0450OgQHfQF6usQTHVT
jGYp8mH8XqRUIM7M8nKLosGIC+4/iRFQRSidgS0to1R4o6F10+mPVuO2MNEmO9KH
ywzrx14/eQYImkTt8QMyOUhOSdHpkOFznTJSu4MIqXSIZ7A3PUPNidUwoYIVPJrK
rrWQWGHU5K3oAwwfp+N/TILJ6pFmt6JeOOmqHjS4hGRbLK/lefSQy3BAuM5Egic7
nb3tTbTQhISpvHd/uDMDXAi/N9puPD5hi2R5nZ226BCRj6cAaGM0HrbmNct4Ki8f
O4fDy1FdTVIVuUcmdDU+PfIkrIEH675dqfm+I/+lxOVSljXhoJsz10OcNtV912Gb
T2jjHhxdS7jZw89ArQJBLgjU6J5Y/E4VzRy6rS+Fth1X1lKxpZMBgnQYj/zR+38q
2sy3adH8H1+ElFBOVYMb24G3KcG3H1qdTXbTMGxC5gdbymkO1uz1y9X/bp27VsNn
h+HvoJtyYNXMFmjU4jy+tLuSRYkf7kVvsGr1xpkq+YETntFSxrdy2kcCp3n5Ergt
x4aB8ICKBrJj279nATljxqqX2cR3oMaSszLkTY7Gz1KyeGxojnq9TT+yxWYCno30
drKOISxmYQ2DcrsRDlv4xakaFloa7jRji5c8vOrGlxQn7SSossN0znCHGe6li0ri
So+p0ck5lV2i9fxoRQxh0awi5VpXTZB8YSG8vpXjeHVoe5BkDoQY2k+ivB2FHyJo
EVBs+kBytJ5aTaz9AlgMfG6GMXlfRlkAhqP48sUtDZBCnnPM9T9Nvm3Zaa5o95iI
OWOVpengC7sWq6/Lp86iJuRVmK15VuN9Y8z7OycyoihG4yLNp844tid9M6ruzIWo
ePfhxsI5gb4BwYw+X/BE9MQAB4qnd0PwwJxmeOCyM6ueUWLMz2IqpvhhnmtV5Ttu
4ADreeNrlE3a/yJdXKFt/z+yJ+EV69B+0j9GhpN4yIPX/Vdy0y14gIMQht46fw3a
ynjxbQfiw9YuRPPFWPHAi9mzOgzM5LPAVMgh1KTDAGsigCpYmNI/vaOzNc+eRowV
mB8GXosTq8wdtbsM4wG8D/WPumE7jkmjkGXtcJio7O6EmvAJcCEywOh9E5BXNeTa
CycBVgVhunsNFqyX5E11UOEFusuMLWHhbggFwKDdL+Z5HXMljnIOU+rNE7oLcDl0
bwEO0ImgYi3fVCUI4ZEYsGg7p0oJH2N7U6N6m//3akroZRcBbwf+72A9WfecO3xN
0UmyYH3J+Rc6TqPMiN6NIH8i+jHYIuCRIyosHOMlIjRuk3Knos205DCo45OzHWz8
KREQdlPw2FqQkTcykk7HzeWE8SKnXOCiul0vnxkeDYr5q7tOQDCKaKQRBdkbi5M2
LUl6s+yaDBZgtYqX1X+6XKhdui7flnrotDRj5koGG/DNp/XMyebWqncuoUDBr3AR
IVG83iC5Lk84sGl91x2fZPYYvKn4W5YMnB2D8c0FgqFXbzGesac8Yar7XL69WHjm
6DOJV7D1DR8jjObhJuJB3iF/h1+nrqrL4u6w0ynvTj/s18t6jw0At236mWBSkWhd
0FpswKklFt4zbn2uc8tYxLnZfDK2ZCeH3E1N3YQw6FWN2pFHGVpOgzufAQNFe66z
7AJNLXahQRRrhQNAu4k0MdU0zwr3ievQRgVoPNv4fWKgbAsKlOy4QShR5el+WywT
8azoAJpnILQ3WGEjEYZ/U6YAL8DcNLUeUBNVMMfXylCiVS02S9hDKE5gK07WkFC5
pqHNCGkJnlpWFMZOLcd/aZHlp7zsWQr8XFZGTaEiDia2qZ9S+cvUyojqL4UKciqg
3YTi+BuE7WR+2/HxaKeo4uEVK1Oii1kC0CuPmhMWwC7QJhfY5hxBa8FgDv1N3sgi
TfPJBHowPo2lH5t0d3lJuH2CXALTOb02KcGkQiWcm+s81oshzVgDZ4Yo4l+klPiA
4oTeQtSuZzPo6RAt3bGO46uhbvKZdAg3dQgCSZEToDWNOCsupFKU+BbnVctpT5DU
ufTGOQbz4tkEgkC98r4vLLTLNGpHG8lAA6MgKGCCUsOURThOe+CdqcCkhg6nbmOt
5fML0S0+hByc0IMU5t+Ty1vti87QzEBLdIkIma8regsNcW0/gP1IDD9nfrfnfOKq
3/ViguN/fYwMvp4rNHvDfAxYHjuCk1qeg0YXQ5NpbMCW2YHCw1/5xIy5jJyt2EKl
HWct8MjmWk+ll1ThAHlat9njiLeRQeEu/gi3Rbnfgqy3XcaaBtIyMkM4dI9dGfoZ
O6rrhfRxMh3Xfyv9G8lC//HfqSxzlUZEcfMbm0DqDcJz3S4BwgBgPttOqtEcJcjx
AJJ79LHZBZDY5Vqb7Ygto25DMmt8vtWanJOopV0EdvWYMmHc6GPksGl1hYRrSR1o
KQFkyO4SCU/xE4j6lMdFGygVTT+aE0Z1JAP96gP+Usy/H5G0hEfmRbUN2P8sUAvr
aP5wa6lZOyKKC/Aya88ry9CQGY9/+ZcRM5DtqFxWtuKYSWNmYy4RO+pxouNoBmaT
pkDbEVs56I9BDecFNeFeYxlUq1rg93MOKqIG+jLK3+wwy9IbAMDwMfdYekHXxXwl
MKJNnFmm81b4n9bjqskZ0Bd/cMwJSV4iPUrf8BtQH6tKj7lJA+ssdsi1+94ljEfY
s+CqMDUQLiHTtj4UsTPUrESDR5OHXOtudXQXfoL2ZCeoEglFBLVrlkmDEiEA3EKg
jU059qMWni33vdT7LGGxy6JFqGs/wBWIMQcoeRlxH+nltITouJspO/41y4c2pLBe
EaEGR2rSsKF4ALkhXMoUmFMqFKUIbVqH/WkH8eAHfc16eZi3AqXOT0LbKxrriEz6
XHQkqhTjB9RElM3MaU2RMoCeBiHOBlg4U2QqJRJ0zcOqCvd+xnV35Su3SO/OXoZH
0bpB8PvGpHho/TiUKszIuPv243FzQf5blk6/mbg00WpHCVpiPmvhXqMs279kpH7S
1aJL8fzFO4voD4yMtQadLzzkkVBrBLbzLFURnZ90aaCXakS16Uq7+ZTN0U0t/6/4
FhssyxYmM61SlrzjHXR3oKiV7N3qq0jwwsSu6Bxt/3Pv5Q1QfPKmqb2ixTW2cijZ
fBJC09L/mbbLAdIUT4UNqjBqfnZANcpTsd5CAbvNISe9ABGcP4J6i5tMmXGw0JOB
eb94LlL4O+dRTh1+rz2LClgR6Ul9PmDj/dH5eHLjyGSWvL6gaKzwq+Y09fgC9TQW
7D5B/qP6BjJwQsA8GVUKa0KaD/n+hedlUnuOTlg6uX1LNUt4vqVxUQcMwx6YNfsH
Xz9ITueFVIGvgwDqVvzJvnjlrUvCBHe2qt6RZPnwZbQs4P+n24pSyXWH66/pgVy/
jfU4hvwG7wF99DHMUTdR5UYCYuOWCHZ1szfLJHhZbNqXjVdW+MSm3YLf+Gw6x0BQ
Pt2wPWxoXEbBlo5H+1n7D2AAS0Ymg+hQuK/PyCcsBvDkDWS8fPQuYotIZu2slvLo
qaEu6R8HhyC31Xt5MwyW64d0freEC7iyDj/MCbJPWdsmL45QPrpWryDRBdBvbTwf
sgV7a/WTmYqFbnRq56EmIB4YPzWIUSpJiEjdvQlZV9PeQNNPHh+Ianjb/EDI21Qc
UdHTEoCgy192+lFn9KwKJzrb1pvOxq19WNxwlnZkl2Cl5KtbvaYT9AJ2MVXnMb5Y
bcQde6oUoGd5iLxLhWjnXKuJs78nTV8l8cTh2A/zhoVc4jQcb09qUeP7rAvB5lm7
MYn/WO0i3cuxd8aNfLnutMfhiO+lEJXrdGEY/EtscJzlRcWWIfPFRZF0wV1JFHGD
je7fY1CCTWZb0/vsU9PchxsJSDVjEvOM6c1eOxq9lCKEbkDV+FDSKpLbylEtQCUB
MFwY81BPR8RTCiYplVkM95vXSCZEa73FbCJfXUv56vT//9XCkBuuDIac8VWOXetp
ySZ0jM2+rg1MSZzXJ1w6ApziRzqDZ0Vm5Xl6gdyk9QvfdjcGxYxcVvdUvur2BUvv
LiyKx4RoGj8LeogIvWKvd/vDns+oiijAZbpBBEgjyKyQmQ2je6aw6amo2qmv74qM
zDv688VCH9XQReBqDuKvgK/97Q9di+si8F2s8Ub0/SruKvyfMKyJMwrN66ok4cXB
6YKsZi/4fyswiFwx8+1jzG59Si/advOA+h/v0FzASPwIygEneDNdo4WjPoxE4LWm
dQi8SMlR3CxpEPXoYDXkYc1MIIoJL8R+Cm6pR1Lp0dZJny3+QGuAJqeghB8E7PXu
49xfP3OQHhId2YqLvF5mV/K436YcArXSk4JNkFD7CujC+fyBn6d+fcVkKiXjytr8
omvJxOaMdmaek8Rl87Hr8vepCIX9eOt3ESQIzlkFYkriZ8So7wwOutd6L1pZCMLJ
hshfFO1e5FF/jpF5pWWpVAw6TE/5It+awzgiZhQuVS/S7EIuyF3y/6vY5mtPtPP6
06niGtRFe6irrhVAA7o3hb2gbCTTdyCLpwlXI9Z4X+ep8xUxTYH/CsmXwA+j+nZi
3pqBYp3CAGPxPmxaH+fm1r7GPImnoJd2xWhagK27mCHk+16zkSHvF028rZcRGLXY
YGmak7Hq1deiroUOruLBM5Boc1Sg806FwvI8jsyRzZZD4lIRq3vk4Sn6Ig4LcQ9A
C/zL9TraFfafF33k1ZXUBlXUJGQJ8Y4cFWdkeHuB5ahAfzkEd/355gu1HejfRKg1
SRFk8GiZFP4rGBCEfiukBD3V1fCaOqPCwlsid+JEljG/9w1g/A7JucIKzpwrpliK
XGau9kxj2OtCCWNPNV302TEOp63X/9JMcyYdq5puSh7Wy1ZjHZ69CA83zYpLuutc
EofPF1y9QAFrNCo5jb2coVjL39ZnOvHcx8eggeejovoi6QsejsPp1fhd8KaD2LYe
TqNj9tJ5A0VAwho7SQMzkPzj/ACAplWAYQ7eDzqM/aTBLjmNPk2fQ0+GywB7Ia7v
nnprha5Paom9P6lUrclKr2U50BEgkUcyj3yw7x3rm1G9g3m0bpdf37qiLRX7BUmg
0e3KbPsQ/xelI3A7ZgZIA5jmLTyH6H7lLMWCc9zwrgiMpGoMky7VEjk4BbijRKQW
orRenooqzknhV4UolIyOPy+edDOQJoN6vnpcrEcnzYzvMbjtOglvwargJKsGNSbp
jttZvbow0FgE5n62jjk/LhTekKYQZHGv6/WTKGW9TK3GlL3WNKPkZ5FD54ehsPlm
ooMnNzNJeE6rPPSEZ1Ojx2/7u9Z5BJtQM14kjkX+eYsV9Mthx4MVnB0KnkQE1Apk
Uv/FMdkDiGnXipbozJ+aelbE89juQr3936viFDQc+5qVjupDULxo0y3DelcTXxRd
eWAGnO/C8iqWmk+Tiqx3BXNSzaQ5S4i71lWwq7KksAVNkdARv4xzgjVa15LAIs3H
LRDXXAfo2Z6dJkeUDNrUIXpGMpwxjTBuU9Z4rsSPSJRuhm9RR7NtT6jDFVJKXH8h
0Ds87xq7AAxIsDj5bFpFv0c4Y/2e3OAPDuTvw8QjDVt3nZC2+jkmgK8ixzVP000f
w23DajMidgyH0AA054hgrTGHVz0DklgmDmwTESbF2O3pq1/6DV5IGk8jg7F/NAZV
OaSBOxym6nftct7uNfDi68QzVly2+ZjWbKnpbJ8piRgfG4Ithe2z7V5h027734ro
4bPwwo1RBp92FbNMtBnqG8uEBp8hedBO1bOXhrFTiUFjKFidTmqYyP67cSMRAb65
RaoQY8yLUbeOujJ4N76GYB1Vn5N/or/Zub7Pj+erASug2JdJAN9hly73H19gX/gq
xuoKf8934r1nJMQl2n7hWqZjQzNISKMMUmPwYZ/QFRYXyfE9iS370TtTdvckbS3c
VSud1Sr93rn4kCDc2MQMM60lW24lMdg3wj4GLBeoKsKYdJWHUhYd4GaDEWQMK/4b
Q0UknbVAwVKFyp8ELzd55mETZxWHEso0+7o5L81Iz8rOlRuSHPsLO76eOVC+Tgb2
o7skeOB1ZuOH8JJVCMvjn9qIz3iguvhYl/0+uhlVrX2aeyx4eES2rqh/JomlMklL
E6Zaju5G7HPieaHBcACv8WBQlEbOpF5j1KfhU7hxRGXocCYJMqh+bcrvkdfsQNxe
okXWa9H0Q88aOPeGyNNrKgtoZvxY3YAdkexVeNFWv7tH4D5WuoJuxy+P2t3Pm0IP
GWGgWnURn9Jr3uhoSOlz9+g9ag33ruYrGSKeQN8EfYDcFKhCVY/t7QO+InDOslKN
bO+UlvEpEhk+GlpEWP7tWTAYpwRMIHg16F47b5yRtehInTOKWdXLlOyjSjw/fCrG
+K08ZYeM1Dr0GRHVXihWeVihP4YK7+55UGfltKGX3ntG0LQiOMhVKewVI2pTK3mX
guUdhOb6hP8eWCVkCeTftQeDUyLOWq1STNR9kyM1BhWdEmBAAbMZhwRplP0M+JRt
tD2HyBOc2WbC4Bbx2PPGcB2u6T3z7izcnxT+aDMrKf4R0OtU7+v2zxzLEXIosN1U
0l5ztGT0JNPw5mygzSsvgoxqXHSFaa+LN6w7IvQUdhU4cjJQ5lF9nZ5c87aFAKQT
xJBI4/U/+6dxA9dh/zIKzg8Xh6SOGDXyu3M5B3Wia4X/wHPH3wDQ8NGBFKRgyn1S
XV/IY6n6ZSrJKdEZJhL2CEE/z2pDTW7h2qgML724hgbjUdZ/9ZZr4dMFW4GlVY6R
0YDh98OhZ/kasoAQy//QekRTBR3lr9AU5tL+ptP9j65h6rtiAM+uIJdQNFbDIysR
gGTkldY0J7SEPFIYyPUMg9TD7eAr19K6a+VxTkO9cfLyFstPZr5rxkVYpGkCf10e
rMT4HNaqACVZVEi6yPdyN+DEJaDXARAJRjg3qOT6q3vQQAKloRCdSA1jxCfmj3L9
a691wzCwbTywQYwb6cpj/q3RzSGKybTUhk9kcx8olxyEBL+8flYofC+bVNSGXK87
3cpeIntvzRE5wVgJaBSMugYX946CyXvk1MwDVvFcDG+ZSJZ5MWDA/Q27O+38rRcn
2kojfE/qwTMlSjt2ZLOZ3b8V3RVrP4RwsNbUC4KMK3KPVbCr9vROsdOyNSKRov9T
lCqsIOmpRqZFvauiHuRN+Wh3ji4TZFfz1yoSIBAkVuVXwMRU6DcpZCGEaaNQEdoN
6qh9U9181paNVpQZ6RkPY3m75F7PZxlHkarhsizuHF3wKgwXPbP7LF57plGErreT
7nVzlD8aod/4s8u/Q7zbi9t3pD4JH3eT0DlJ/bCVxT8m607aFlI4gzUDZxIqVWWr
JNMCEp3+ef/4cyChj0SBDt04ehuc5JZkE8xZ75dx1ff0NKLEHeA//xVwi9SZrElj
RJ28IlYF5Vgm4QNje/nw/vq0RknDEdVnnttF6gANg44RqPloedgX2Q8SB0LuQlVD
bo2EOLYcSNLeIjTTsl0QwsKRk8viw1e7SvSGE3ChNmgQnX+SQEK6WLbw06P/0chY
vfAUt7L8vGsnvgKsuRiHQAwqQUQBI4FEUAa/YRxIN9bSJAv5juIhtbb7Y/5KRuVZ
JunICPGs3OjReCRDbLBV9KydWFYiNm3CiuWFFQPoz1Oxdri0N/j74DHfjvk+3y4K
yNSi3mZMsy/0hxCZDZjE31e2OEeLL+7PVyDb2D4jKAvmmnR5OxOyq+B51+0Ztfs9
EVdLsmeC1EFajf5onTH1QP0v/uKH2mAYfniREyCaTKscI30eNjrg2uEMFzwdNpTh
U06UBaeK6eNhtjpqEDIpbzrAExlK5vXLmGqQs354I84jujafOvP+M2El+6qhCMTu
yHgIv/IyuwcRLRVdSpI4Op56pJAF0tYBzjyXMl6w+oC3yong7rFhG0UT7XFEmGPx
8htrj3OjE9Bqm/NumaDGfLipKaWY83LpI3H26k/r1UuCMRBDedmqRrUiWE/2MkUK
mk46ZDbhYotuNHDQYMi6d6bZdAAwTU6vp+4+5rWwhzMptwaUhnA8q57vqySCmjTT
YhyFrGyQzykWTyd6WMHHk4tDBu1VBVO9wPhDEjtuP9UPBdECu5ER9XAiQSfgzwLX
rFVq0qimMgFOU7p+Uojzs0wNr8edRSVL9lxgWN3k9ADfIMKeFwlqewSLFKKyMHtp
v7eFIHAUTCZfGqMfwB9t+1EbGVRrQt5qQX94r3yWAw8YHxUogFf6IvHSm/UTb+HO
mf5GyJsPiEjaaVv1LHyk/SWY6jQK5cwTBO67RJ/xk1sogB5Xfks9deSJHV/mlSNT
tpYDSGL3ULm4IUI40yF8FghvcP+WSbl2YucjZnsej04SLo/pEaxHIlZKGR9rnggq
lO5VuTnSQAPG8JUQziZTeVYJ3gG2Vgk2hloTAY7mVFGf4D/F6JRpRM3UfUYx+1zl
JMa6RrU7IGzOUza9D1u54Yt3sVX8qeA1fLxlvSPd9HlJRBhREZHJEOEWa1jpLUBy
sPqQNALzabbta4jqv6Q9dniKBBpkrcInU3pZs/b5b6AsrbmTZNre8AMm1+8jFOk8
WWrkreX8H4QfmFs8Q6u9cpdHE4iJyADUUFgyZI9yuy8IgpvWFuv0k9maH0psq1mK
1r+kokYQM6MFbXtR5nzmPgf1bzwVHqlEKjbIYvm4tUfeqcnRaHVuY+tIZ8MEqwLb
hnnUo45r9W4afUENgjECvzkMOaoGu28ZZ1F4iB6/Tw9ZEM9aYCsf96NgRRZidLTA
4uH/YIc86xwZgzQM6gt4r2ljLzCv9rYUX7tzxyDxB5Y/nwi8zyEQ5ukGbl2wY2oE
+j81cVospvz5FPaltve3rBWgq4c7u+fnogjRw7XZFLQvfiXFgMexGO9lfHQ9AJmi
orrZDtmQmNKtcKPMf8TpRW69Kt/+CocyZgCNjPgIQqHX7E+QSmsKAcvNYza/dmR3
HPPDt/2M52RC/bOgtTuoa1zWsXLsEkEHL2mt/s0QqMpIhiq3LvMf7iWx85+PIKIo
F6uRAmCZHoL8VIRAL11V4a6qlzDmJGFyvEFnWV5YgnRJ5EELwcLJRrR2d5YQuTEG
o2A6KEfrWHFyayP3Z+2K8GOigCvvKmg2BUrAfG1xfG8SbN5V3I1a41rBZlo80Z2T
7MiU5h34I6mm4UHK2NBUbx3EGMiVzC/i4WQ1sJSHunonuz4BvvlkAGjpK4Fwb0Re
bSdauX+ny0H9ICviC5mdBu2GLONm3PlN/kAiTPxWgBB561M9T6Tn3iNp+onE08HB
c9gjkZFZGQfOVId6GG9YOEDlVtB7Y3MGFwoytB4YP3quPglD8WfL7mMEHj+pOFWW
NDu2cjIoSlwXjlKholU2xLLkWljs0bltuOgG4e3hZ/u1d0uEgS92Ti8RoxaEIlAE
YFxXCwcQ9CYd7qJywmdqlh5e0/Ko1X3DPyVlHDbUaJSb7j7WycFSRm95aYYwj4GG
rFGi3z/BR/LhvMsu1LWW900oTgE/80jvqiy+74zySncl7fadSeWa7HVvFlccgHdH
UMxZrgqxCL5S8OFqdaYuKR7BGnrJrETtLczLC9HiJfIZlR7q+5WN/E/P6iSBm5PE
lwaiKWn3sPbXok7omHwqI0TUai/zW1jUD9TWeoVtgGYmhVwTg/0j8IQac+ag2eCJ
6X4lmlJ16AB0+93ee+WLc49oEC8qsfuWY+5+smXhHoOk0YgUIGaZBqugYYHVn+tj
DSFDrWLUoZuV9XctD+Lc5PXadqvdW6yyxoNjc2xenKsYYwPew+weHxoRyJRXJI4k
4SUxeiOA7/No7wMm+ObuzUgMpddbQpR20TgGCKCSthdckfWU0ezd5EgXCHEdxAqG
GtbZK4TBDW8wjJgBv4iePX/RxrCdz9g2tCndTlxRKHoI4DjHX0Azg+dXLs9Kfpfv
Dzlfg3/2HP4kMKgzS6smt64UdkdE4lGRKIKm9KqlbtfIdB65TTctB2DSto1J4NZl
onvetocEvUzWe441yG+PkY+AbSdlgJN8yupQBn8Q4MovoMqRfWv931J7lytRpd2U
56z0j7Yt0xm8QGBGxADGa33fEMAmphf8hBnxcOu4EWIPToFLZijKsSLit2KvhxTY
Z13HJbo/8hgvKBAR8wosJ2+uFssWOpKsFdCs/C9Uh5R4sSMgE+36E5xmelB5hqo/
Oi3IQCSAwLGsgxUoxWPd6A72jIOQNwJBu/rkk2hnfI2fSX0HcDeueGNDfYHFUs0U
U+rjN8K6M5HOBFYr25CWmpYODwHkwtgXgocqG6Z4p8mqps7ySw25p8invgdB0tG/
w51wZXbkcq7ek2CxpDLFOgWOOBdOjMC7RrJ/Sfhd3IU7cxJJqWOiF4H593tqVcM5
5lNNeHogEscNE2sRFC/YTq7fQckZ0qOr4fpsqLY0Jk6r29YMuj2T8FYXRF/jVU9p
1vr/x7taUaeQbOFyLx8c7p6WStayjHdA6bZmCa4ZZhT53xviMXXEyYJrPT6FohTw
6kGV93yKLfeSvAnhTTjIuPQKS7uNjsCysUWbDYQ2Lf/z/7HjmZHjCq80CeCnALmz
3pXAbDu0GlPDI0MESWjfBCJwc+tCJ8ruqSzGL7aVyxJozfh8CU8b0VO4eQ8PU5mE
Fz6Lw3fEF0wtcMwMhrALJYpWUdtmMOaYMkG/J8LuSkOR4ghHh2mxWzO7iqjSitwy
wAnf1mHZsD5TrZhIIl3SM59mlXjB3TCrTjLjZEE7AwXiSa0pmetfWDZV1mUssyK7
dniw9GCWpm7b/ifk72P/JVGEBnVPY2UCei2oW7GTpUbe0MinWGGRpYG41ED9r9Mr
NoppsJzCX9QPIJ/nop94IO4/CnILFMqVCV7+ZdtbIolv6Jrs2qZmrJRVHTX07lQU
6tJ2x2sABNHIJqlwlyCGNxiFpLlj17bUsYRumamU8+9Gjk8RnYrxr7WytxncLlSF
TlUEqcRb4AThKxeuF8brtqRA211VG8VxvNqlXeVqyNhNTlht4/PkOxNK4aao8kfl
7AYWlKhU70pmgF06fNR4juCf/ox5ViORdSJdNyyKNA7YA6z3oCWj6Jjg7Oj9gE1W
xuxXraqOOZaiHQ9CrkBvk8GmKYL18rfyzxIi72lpXQt1FQUcBlLA8xKfzKEZd5Nc
6jMEV/32EueOLqhN0B3VLJtYLMJFU13Ir913+b1rouNc98GjheRubxLKjSQjxm1M
0Xx/nbaFDbyqyFgCnFbu//BYGzeVn8MesFAvGHMADWFWgq8bBMnTrT8rXUzfBv5q
C9GDotRh61e6HtcYLL0F5p0FgyDAFYFAeWslj1O2xSqlpGLiB9KfGRsSezqPp7+l
JhKPCcrB6OdkUuAg/mfknEpNsxdoii6rNT79Xe6rI5nQiYwZoWst9/bLH7VWCGln
IgH0z4/ofvwBGLTY9p6206sgCW4IZG2SJfHToIAJsy2Taz9QT3cl7ugNQXghMD1U
8R+FyD/O+Qsv/WFlvZX7VmTXl8OhndkxXBZi85/eICOI/Ojb3bXCNcTcgf6h/C+O
ZQVITfatrAiCLRrwED7hEHG/8n4A4tWq1JkRm7Hp2ygzteVWcH/Ht0fvEPOU3JTC
U0AWuRQXDnu7DljkA7Wf5CmypdaAFNYtvS+KNiUahAum1lkS4b0AN99ja7KaS0c8
okHPorkUNHIqhER4Mef1T+FDKgI07b4dcceaSWrHx4yjB5mh9ZUgolybKYeHgcmU
lh/k2ccMPEQQ9x8H/Fz8oGY1sreVLicYNpW/lYObYvFCoPzmxGqMCegaPHiCXBq9
Hd0iFntCCxyYebGDWtPxzczX1aiHVmUiYBEH1nfzOpzy6MPGoFxUIivtX0ILN5VY
qaEIbAMTvUJi2iGZ+mT6ROtVs02TxF8L1q7VbLGZGAIZw27VrkyFeBj89348lGMZ
Q4x0bw66Vw/rQojJoBBs/pRtWjIAt6ZANOdcNru23XtnsROOCP4I40hjy+jH6R0f
96HXAsN9K/DxI/TK3xKdJ2hHjzHMrLZOKfFwUUJ0kK34uzaQuq+uG7MdRKE2RTGS
zkn/g3Xs5rJKfB+sUFayUJPHmgpkRLoGjjkgVuassazNKJVIegSytund8XvQ5gTu
muHBH1n+Rmv7qy2X4jZh5PLCNIEoNUCmFFwY7ZuF588Q7S+AX8ltkHjo4SywocgL
b2zYIeUW88gSGlzRXM9mtJDhN93XlDGNu9ALPWmjAMcckDGL57SHo63A/GQYxBmJ
t2lC1kLALgMy+FnvedkBhwN3QxgLbBaGwlzRbUgvXXeqnZpiE84pTKNieWnr0nKs
v/Nvpfa8zvt8QmI5qPccBTUdefY0AwWN0ExiKMfyy1su+yG67ji9wnGLXZfMK5zh
xAYBgvWT1gTs0tgA0Wbl9drRMJZK4gcto7x9qq7zkddzjh35gFk03hzXGmzIjKyq
jNBZqpdtYcCB05lLGinAiBHTUBbcJAZzAwPbcBgbjr9gc8VmIJBgqZsmXAaEJyRf
DYkhaK+AKkilxsM4deFiaA4wX4wAQEMBHenE5a8bk0lNjRqRdbwM8vl12V6o4Oww
JhxgYbw4zEr48uYU/3kKVQznfkTlWlsm9ADF/0JjzN81DJQdsr+4FYhuclno+dIT
tCK+ecL1BmmUFQJu7hn8+pF3Ioa2eAhcnX7Fj0f5KvMW8fwjBCb4w5NHxVSgdpcO
uEDekFyE7SJus4sm01DjgS9OkH+H4/dCPn6npCKTqVbbNlB+zefr+YOj6xqbLDol
N02ZbvMfYMQ5lDBGtH0t9AQxf5x27Gv38i1i2e+HvRJe40K9jAFHYg8W1FAvEkNN
np6eGVBO8/QRveTPtJuINAqO0lHURU/57XEFgVflmTej9biTxwOodVQut2QcemXv
IE/zgX8c7/hHsj/VdPC5b3d3p64qrhGpTNPb/ifqfSCq+T5XWH/yY2YXURETFYWt
JKYBMC44kmopaCkc8quhJdUCZEPA4g0guZFw165PSJZ+FI/bJwwOrcfEa4t4hX4u
jPzFuHW0U2T0bw4JugXx877DaqhvSmXQ0HjZRojgzKuNK/xgbgxYE/Y3/weoDLNo
J1seI+WWl1AmeNsfSBLDaohKpUSYVD8wht/yoHZa7txtawgH4VDVAYe28CugSdDZ
VrLkjCKaiJOHgAK2njK90evj8/yZHLeueKtf5JWYLymZRSwo/cYCYlT2P5p2PnT7
C6cQ5j08pNLJA/hWRYjLQtyMYl4nUdQA+LeEuAhFSk8vLSYN2w3drWs3XCYZay4N
KONDFxyqwu5ysmZ8Grk7Cx45M2rNy2spvcuVL90VpC6MiKwpaOYrNvtQPY94gM90
1xAEWhZsEwoaCAoV3ELmzYo67pKm+h/glwmB2kusJSKKV3b+vwaqoC5kurvqNA8R
vvzprsiT7XwcwncSid3vN88aX5suTtode4IbBq9EiQ6zAzf1SB5bliWo1GhlH0mi
wN23t46EStcPu8hXupeMw2yhTWK1C68VflHOs7m+QA/tI9UyDep/oC09D0IBA68l
TNYScRDe0JYNUafpCE7knEeH+6zVol430rA8x3Vj7/fUomljFiZF8WzuSjb19ber
jFofqaAwlu0BCMvzP7j7HLQmEV1/ylaemFoKACIT0yO3o2VB1oL5scUb8Vds+N8z
4FsAKaMNuhZbgvpgLX0xv9kb6ejthKC5nLUIMmYLFfuSaOrz0fyHi0p3U8T1ZdQg
bIRzHL9Hoxr/a0qzqZTbXrSVVHsmTnOQck369rnXctfIUKzLnOXvk3fV6/Bjq7/8
mBLO8zI4neWbB1saFgv3k/2QmHJYmHI97CvWreajcCCybTEV/5eqII8Od1pPjQxG
QrhaDiuXecsXbTBKT1CJ1RQO9GGeEo+j3bdo2gGcFVVw3NtW+16GBLHIecSP5nkk
lmv6mCg1GM41GfhC0LwSybPSxufkCxy/yKES6LTJv/yEupGlm5XGercG8e3lAZXu
ZtvdY4ylD5eAfBLADYl4/c9ovy69LTv2sOL/U16X8Nf+gEyvFZjY1AoWHNFGnAdu
a9bJolMYTxETWK2SZ9CHAgE7ufgK9RvQJEMpc6R1kwREdJ++Iats2ZHdLfxL/VGY
/161NaGOXObbINPPlQZWUxBDb8tzI/UW2ujtR2UqFsMnpmyLqQOMtlJdGCwzbRfv
WmcZcEsaKBPKN4LSCHPyjjDJsJfICPl3G7lRK/QdKEl/tP4Paxe5bWQM4qxEhzrZ
ytQ5pvuP6zkUQhoXCSo8JLZjY88OTQ2IRMDrZkSwvK5YJajztMO3dphyEmm42RdQ
rNbNJx3gaLS3nK4UWgBXgoJOcn/8c1HRQWNc0aW5e0I2MvtEv0izc3382mY9aE6w
6wMd1TEwN2/t5KM3NcvRutCqG6eU/Xh2RPtEusSlPujRLA4B1VMhG4DRWyiGlnKx
LpkhLv49ekibNE+J+CT/H/H4kj2RObv81ruTYAV/CHhvYRfhMULQTqE0d0zwvX46
AhmtDSIDCgS0umcKpiEYgb++dwAZB5OmcbIjo+N4gkkC2kXdeOoT56uLbHc30pXZ
WOh24wOPsMRrhZxr3wD5ZNNThqHNzJrVj/aMzRziIU1n+LzF+EJ4NEEVQHIXcfi1
KZJhIa6bC/JNf+QR6APgJNFa6AbAfhoOmrcf8VFWZaRv74fFD5sVutJL/+FPYFom
t/11lAgvvdPXV1W4tO21WZIEQ+75FNUP7tFGGGvA4qszNF4Ap0FHYD0bGYAP2U1z
g7IqBtfe/8jv4imdPRyzOUcW0ABTM9LsXOaxvY9M7rvXXt+F7HQkrHdY9TmLY8mv
SNAlfng8b+vlob8d67KxnZJki9x8JRqqB8p5iz650VV4jY41/LmJ7MgZOqH0bcm5
tHmyFv1IMH1Ycl4z80nRx+JrBwKZudN+o3x+0XHjRdxb+odtaveCT86KsBclSf7k
QvCKe4g8428b0y63MpqSTHHgFeEfUSGO8T3JJNoak8KiNUBumCcYa1CSem9JbiWH
SLk//ecGcD7XIvHcM1b8ZLWuAz8SAKZYztsDoJpkiXkg+jCdw8qMkcO7TuQdWfA3
u/lniW6QH7As2AIlxRJ45lQV0Xe9sjCcd3zCVad8/oq4jHaAUOx/1lOcAzt3pjlF
mW5k4uPyNC0goS4Eg+tH/pNt6skKOE8sjZhJZKHovuqYxEbmCgvQDegQuiI43Tyq
5oN7mfoaeFEkycRDqeZnWe2cx4in8MOLV9nG39lGCPkHQ2LSBOFD3789sa2lJXMi
bdkZPZWne+kplFdXLIfecMOKK1a23fVqbEEpobJ8KFc9cY1x1RGm6rzdCn99itYf
+1+xFcQWq9q+8TeptJ03EKBPXx81PmlYu5SX93EMzvb8Foi+wOq6d6Q2OVTTqMb6
1XMB44R7cuCD0O82p1FCNi/jhIAHTAHGXi30t7EVotc0sJE6YGLRkG6UtrK93DAS
xzGBrj4FpkGFZSB+P6EzkuoY2qSnkh6L6RSttuHtsIDQiWCZ7To4Sz0cz7m37SCJ
yb3sVDZ8Q0d8uP/P/fKj+OjTGOqtc8G2iVGYUie9VabNqNoaC4if4yJtgueYFP65
H9WPM2EUrWyVXe3FUln/Qyd1Ds94ox/9RtXNH3rOG6RhD7zSLzRF4d84Dk+MgMFS
ptcLbGm+qxeqTcprS0bnCnAxpIcOxmdPRdMYrvIM1fddMCi3hoVl7oWYGHVKlioS
wF6bCpzPfZT3sj8eM/y1TakeoPn9N27MQICuHgopVh1nasShM//0AzUfZmTqp/if
381vPWZzpkIszCspFzr6JzLmE/IQEPhukDsktAdvmgijsZonOyn1aC++4ncTtvFZ
0IJtnfY+rXObsG1srvv2pYejPkmhXFp4us3JE/a05jMhkitDmAWOMF3JDQqN0iIr
FLbYX8yfImmvYikyYTzfVHMAqBozRytHpR3i+Om4nEeXgDJequYr0BPWjWvD/OS0
QU4lmMz79EX3zgo6eBdnhmF9fcy3s2yPkGuQeL1KLXK3BKWSlCD5VNV3LQPVnXni
UYwO2jSdBeHf3mxQf0/JslBsiP0WwgdeeT0PGs2ELsbHs+GlPlxtqo0bIOht2LrZ
oZj9ZDb3s1dwRB8S5een7jASiUIF+rfuh/MadUI+meW88wc63GLNWN9nlLdb1m8t
78fCUZyR0ChdZzUKzdNot8921pfzdESkm10H9A2DRcybt638ktHijpTMcR7HrYM6
CNKIbVV2NWCyXeCC27XGzd6/brZcr89GNP6AJgB1Eljezpkz2LQXIjA2IN2yrDXV
cEStY8HlLYEuW6EaLSonghXFF6x1OyqUqWv6EBKUiT2g0SqfqnscVs7v1eQBt40n
TtJ7VpbHCMkibi0aCw5+Fjp/tSMSt6qI2risItXPdKsN1rEZyd/y3s1xCZelJ+CH
n9LvDgxC4fqJMDjVYZltEs3QXPaMWkCBCbFWtmfAUgfDArnnYP5OzsXl9rutDQq+
dGi20PPT+e48jqhfTx6K/tGAsyEf65EDHEuJb5WalMpK+LsNNlEFz7h4OnaeyPS6
U+XAn9xK1yXi1voQBfzfQ7DzkuxrSZ3XmERUbMdw7MI28i3d8Ge7mHhymXJVjBpw
pIh2hKSPc9C1RErpJahlNzdhMxlnssFIVL6fomPDiyS71cpmvoDBjiBGYUUAwJBq
qf+/h8UIOkX9X5p62cPvBModVFPv8sVyE7ZRvYw/SAly42sNItj2mnvkEZNf+E3l
JvEUp5TzFvDYSCbIgD4URx1SI825JAhrIkXw/xmTJ6zHHRDeQsZOBLUbvY8YPMUg
jUuMS5mJ5NJER6cxpzaKN0s6w/r85qBrcY3VrSWXL2r55opY6EFnj7cLE23911WQ
loE+xtwVrfQGlfPWzgURPyPTOQbxUiUW5PnGexP2t/JNYVXArrguwCYI8tKS4OiO
FUDxNhPGexC1/v3SEK1o1ijav/nXKptk/FA7qFBeIV2EbKBVmFmxYGaflf8BQeVw
an+G2Ew+KwUXYcxt3UvQRmsBLWhG+tTZQw0nKYZuQkO1ZHKCMsTuQWuP8nt4XliU
OMLdYXwiB8/Lkgamv4im+uB2NSK0BpfWah6FYF0TVt49FDexeqkzRSZBWY2X5+fQ
zhK0XuWhgiwzC58ytcrXSITCMyXQXEa1uw6P5FXBhmAv2LVrQOmS/0oxOSlNrrJY
xoBRmzO27Jh9dbhoROm2h8SZm0atN46gXfh03wwI1DNeikV6IxYTsCdMs4pyyICX
bSJ8k4qePtAkxZn5kdZuBy8xwjBMYTPlg+iz0gC1cC9YUcYfG5DroFxg8V6s+OCR
lycGx3moIETVXyke+aWUcpecW0NtvtJa9OZbC6k0p/hjQbwUgD8ip9Q1KaH8UaHp
ms3pltZuRMKC9UlUfi6iRL5KedMLUhqmE8hUK6H5SUUQtOdYuoFD0ehwm1WUJT5o
/YM0aUgy+AU7BvfLxwWgx6giFVvAvjhl+wwW0FkDx7ncJU3ixPlm6bYAfDhZWfgO
P84GrH416sNjU+wjCdArQKS4glhUyyJ/eFJENxWPM/+6e0kP319f8ctT4oJhkAaG
qtO8TR2HMem5gkGJswisr7cFTEmzq3nUuw8iQ8GD4u1tnw5vzkzBWP1NWmh05cWU
k0JcW5jXhudUvUy3FIVv0s1wPiuSc3I9Nq9tdARZNb4P8Ub3PVTkQ7fKTPN5Cn+G
Z7x9SL2W1CPKbGaas48cwdzM7kTA0ASQ7e+p64xrpmAf4wEz9fcGc33zwhzD+c9P
BE2OZ72+UlgCfYns8ZN6sdaW87GQEpDqoee0eIrV0NAYOnqgywuTnNhuoFPuZDpm
qQkjNpbSnsB5fys1uTmew0BC79IA5umqh85nnJGC5AumvwSDUDdzEdgaZ2A5K894
4yVA0gt1odXOV3B/hOnBwInAj+oxZpFgyuhGmYO6W+IJeB96BxkHbv0xl61nl+9m
yXYD5dbqd5q8ZFtniTc6Tsiv2mhL35ko/OkENQQzuTEdwj2Id38GDeQe4cyoomGh
TvXd4FPJ0UOdT0ziHOKUtQsCs/RVYdIJQLrvgHUVUDz3BPdamNdRa1nfjI6zVhL5
k/SmF1XUGk936kowMEoOlaxKJI12bjVMD2UmENqu00cGzFBjONPYyu5S6Dh3jdQ7
K+yoCj9yQ11yks0tunGNHHzrGYR6rQP+Ttdn8Al1X46dtipiZDflWKhQs3dhpD47
YVv5DL6X4P+HfDDl7XpsKAC3/BEjHL/inDdXSvG5GHp3GVOMTiEvZXshmwd+sJ27
lxN9Sv19v1pjpJYWs0ZhM6Q6iE2f8Hta2qBaPmJSQOpZxeX0eADUjWMK4zmKnQqI
PrNElhZ9qw/nOU2PqjwnQ9nw5TKkN5cRW/R7R0RvmjGrKoaYT5Q/B1qsNZDk3Sin
tInycm7MlmSfjk/qyCZo7ZOuj3/aEYd1ucPcmSfkV+66myWGQuHW3u4TtIq7G3Ja
xHBYiS+fNY5HP6540p5a3vZP/QDsqmZI6hNOQNxfW6fNgG3VNbsS8kCXG8EW+Tgg
pUgfPKUudHw7P6++rTPqozx8eXsUgbCHCr+9bWPwQIAmev2oQnyYWUjkVEiOph56
+1eVG6sgNLvmLgSwc/Sn2cWDcd1tMvv+JUiGvC4ojgu8rKh24TuhoGyzd5xAxmRh
gi1vTE7VeJRxHufVjLBuy7QN/yZYvjPbQ2yRib4/gyNUu7dALggQA+8O6hNxOc7M
imUq7ywxANDcd9eSwwF56/52Udw325oSRuWNodOugqDkL/W4UtiHsVR6iIjzNGtD
O2KlZ86qFfmJHZ61MEZi8zWlPh+W/q0Tjbr7+N5tpSqdQ0YvAG0fCDS3RUvTrgoG
JJdon6Jk9uK0CndJDCyd5xqccaLR0MZf67N+v2R1mTJ6KnYZdKvIVrid8bN5yTsj
R10jXxbJm/bD975Lgqp8rXtGQ8Cq8uwwp5TzQ/s3+SpZOsvEAHRIfeJu5zP5D0hv
gvyxLE6juzT7uydl8g2kgjHbCR5cEfed0zIzmVG+/wOmwwXkHhvWyfwe9saZoX0i
SqwyWpaRWxfAbtDyAHcOl7CbM+5S5ehjspaI0GnDSH3omOlXFiUzvyDt5tUdFoWN
duRXshcKBi+QjRFGh/JdgcOZ4j/V46tir7z+CFjJBhT3/9nk0SUEbGsE3UVNuAND
8ym9mGjbxyxhw6SMA6OIFljWkZxfo0Us9G/NBMK1g2Ka4tIxBaBvcoUqJcQpczli
ceNoGp0GNWXmuyy6zmKKET4syMEnUJzIY+Nnar+yLJjUIMtE2KmyeEUEGjdbHj5h
0NVMJYJwLFGYDksR/iIXwNlh/MqpV9jAPFNHG58A4kIIFQ+mbYyRzIYcFO1c45rV
p5MwBSei51AnOt/VZ79RgcxBb8vWmUV7Z9p2IqXx1SsYRpsc13OfpQC76hjMxpDZ
yiXxxcyTojtU6d1DMn++k2yziH/q2ykrJqhemttaDZ6K5im++OW7DOC+qNTaiNYn
PlaC+vOu/qwQKy/xsxpmnK8TjY85iK9qcMD1RX0yECJDhXAYEdjW+rzaxSChS+ma
Wof+y/0PqtGWxUtlLW+hLNMLS5vu79eBc2A0K2tsNJWPl5fXy+CwPVuxB42KlW9K
d+tUPiEtkvtIZWefU8mVPcAse4EFAlE4tTfM+tdjvm3N3A2PkyZYZHoLb8Ii0AwR
JznHBguy7Qom8K+nuBNzAH10R+ECnbk8iOZ5DHlS+7zJivhNaxYyNZ/+xazmkn4+
wMJ6OFtyQtV43KdCA8Gb8juDGBQQg23MDKHYduZ5afh1SpQz/6qRfWN162fmDOtD
bEHpcZrfOpQ3YqJle2T3ATnJUbvSkbIHECrMVqDSVBVm5yP2oJIz2DnYxB2i5tmE
SrCU9MZvwQYOlc1W3pxNipGrGGSrAwYtPc1L1PdGJ0Mh+HdWfyxEGQdbsPPXxOpG
6jU683k9kx4GzEozt0oRqqxP9Cv8k+5J+KSHp49gtomhZJKZxUlmGfSJ7wdmQT3t
/UhwDKSzip722gj0pqgBKHk0Gl+kuzWoMZ9ZMRE+eu6HCymPVbjo9w0fAMpBkmAg
FPbO3VeUr3a1IAD+lUqF1vcPly7thWq+YU2aq+6He30n5U+vZVFl/ET+lu1vyr0k
IuGkSctyxMNX9i20tf4UpImd6/lRWJsrlV9IytkgDtjBJGeVNs6otTJkiueHKN3D
m9G0o8APO1iVCnzJ4+GiPeSz+r1PsLbh8D0uGoxJ2f4NMgW6h2+MjJzhgO2j8s1Z
AfjLN3JiLsdz8Y2JpUc32fNyxVvtuaBEtKDI1+2SzUpuvdU7JKYFioGuvyZkyZkd
DDBW8ynj0AuuIol4649kBUnTYoBBqDzipeym5JKQ4KnMT3idrv1Z3kOB6CiuNrGj
sOVTKN4qU424kOko7U6LXxFoI6nrTL5W5OPcXmJ0uzoD9+m5mP0evpJX9HFdU2ft
pikNVRY6m3zfHA84L7vjadl9sB6ieFe5RcRPMzlavx2HI/AM0F+3TxBHOegx/XGF
4njjh/HtoYQpzHvqIw713Nu5qKCHr3MiN/m0naDvmAXQDEuFZ6E+gJbRArhB8hRH
3b4+kky4Fkn6jJdxKE0ERAkb++XPPE9DoRl1+jtf8B4Sk3PJl1+3DABIpP6zKy8T
/iIIWcGjT29rdd4cuzbhHmtdRs63pjYFUr5EF5HMFYzmnPqGum1sdiVcJhtoGX+g
nFjYUWz77YeyMm5lM/jzdQIaf/EfIhnnWLwmmN8foea8vNmZs0+giw/mUPn/39vq
a9fGBlt8GtFRJyAyzK276fHs+nbHEvPLYM0u6U1loW3LdlU7GFUTw9gb4zEXevIs
K1/0t+IWscYSAjn/miTy0tSxeYz/ucPbBzVyB6GHMtE4xICOZ2pg3zRWrz8Alx51
71hTbS9YTjetMKnpV7tVTifTMJtIqsTWBi/0z4KRZVR3Nu+Yhsc6kTpKzsP5J/8/
ef6jA0twxw8Unafc8QOeWRCmM3+pMJXL4gwjDdKgFzk8M1g14fyttgw7slhtbP5O
JMGjuhXExSQOwSXPrwQEUydCMgprRaxVWxu4ISPr/qO4ivtLpveGz6GPBWaYWeSv
cWlelLLwPfl55CMH/AVaG9ro4y+QlQDUk4WLBKQB7ujgaD0WJw5HeHKVCd/421YB
Sq54mLMEpZSbWfp5P8T3eD8f1vZifyEtPE5Vw/ondQ2jUGRKUesi5SepstgMby3s
3n7VzI4FHJSkuGFZ/TgS3hYwXE6DyAF+6/Q3Ohb1rcNdCQubzuwTPp+koA6XGdUG
Tu8pCPNYOcfMeGZ1P6CdAOfS2GPqXOYTHiQV+ob5pnXhqoky9UuSz0JY+OOVIWa9
W3deLAONWfXd2zv7TFt6JFsU6KWQ8lqQxLpy7vGtk8E9lL/q6XzIFPhGbN+1J7Az
GbB2B5g1mFEV8gTVlkjCXvXm4LDE3YZBBMbSWccbyxsIz8RWGlqKN1PsJ1BlsgiB
W6tN6A6Vvk9eJLGVzzpVoGDmQnl4fxmw4yNXZ5wB9MdQtcYuJPfLGhFyRYUVmMoo
bt+qq1sao11ACNLlh103sO4zXE7DWUks85uOZoZihxcoF+/RqPadutPZXiF8tgbW
5FbXRkNU7ZdxWCvohb6Swpty1WZhrGpgnCco5kIix+KVyzCR9EPaYZfYhDPzjdyH
hnHB1my6PtVx7sMSHgg5v6ysvvLIYTgiFVt27r+4SoSPWA47VrhpzTloKK/VDXF5
KcHRcbIalCgQvv7h8PDmF+4VeyJSZ4CjwCFEbYd2UDMkgBqph09N2lRVksryPUrw
n4u2lc/UxtHwiDWPvpMN1I0ruGcPnwzf8p1NhMYqS2xDZSfUyaZ/spL4eoCd1TCs
zncTa+5Wer9R9MYd2+ZF4AIqKWbEQX496VG0Qv2eERKO6m5p4DthuWsYfkbGz3xS
68nxhD1NfxPC4Asm7zMA8OlmFhSyKyltWidpZVY6RTrh7y76cWMtRi+IrCkZ6/4h
COKwqeKv+SkqEc1pKU00ss97duIPNvCRZMWvN8XlJhrlNQ+UbJ0GlLiaSmfFTITd
hW5oacXXHC9Fnl1XfINOE3qD2wnlz0aDrAmAyX1wukHrRHTVu+Jdi0j8hFgCPOq+
9ZgIOoIBZ7HEC/775Y2T+U/357S3G6lMWgO//EKz0mMWMd3zI4cmPoUdkQsIvLWf
AHbxEvdNfNWviOlf613xhfgzjF3iLyDQfh6MaoriJgM5NsQNS9Zq+zg30zHpUHqt
atzwv56IA659NS7f/1fpVykUyPVg9cYobv8jINgb9AgNI1QPM7+ZGNlzJb7PcJHB
On0efobgNTsz5Fp3ZgyAaerJlrm87lYlNj2LZS84nXiG6NPw7TrCJ19iTdfay8lT
0gNQ7p90rvOYFM86NJa3GeTEE8jV/ZqMrlZIs1/ykDA8vuwSXF52T1eRTNbYZqC/
u9bw1tu8GMDdXpIw/JLLU/5myLtaVvRx7LGTc7zEZwV44UJ2U8+Sxw7rIV7kZrtr
anSHQt1t5SihVG/LIbh2z5UrwdC9TDF5jOgKXBlIt9ZlwyDRcEMmX03GtbfTc4TF
SRGTpvnXPzjHWtEi90inkkY/jNSM136vq3wgyaTkRP9O7SD12uNeq+xTsI7aqUlO
ubEINvKtJjjoZ+BzVFgIZsx3hXoBzlZg2b9a1glAuoTnAAxCZfAu/2H9pgEgAkK/
hNt6fKtvscnskddhe3Sr0Ft+xWkhwYAZHz35n1nqpeIWVw6PQU0DGq+pqhTPfoC1
8o+ShCqMfYXBjjhAHiigd08P2rhN/Dq3xkXvvh9VNkvzm9sx2xKLbFR6m7Wy/1HL
PwJq4tH3G2fLML0WLvW13DSE0BdJX0F+DtyggL3o8u1TNyahXQG/6HsOJJIpwTQU
OA9F/wKJ+FJ4tvewJrS5trK0BBaLRQFhyobaox7x5MAp51XYArPTC3pY44ZuzHe8
Uy0oKIY0cX+FOtE7kRcPkgy01UEnNLpzo9e8MVZWYeMIBJXc4dxH0Cy+5AD9POez
SxWgiitMzIw8xgPHnBkirssV0R3dxsAJWYaorvmnkYd0v6M8kY8bAGThK5nVbgSk
BDBkluYXyTZ4osC+p919QcC8DLDAHUlcWjARz3DwGoF8CSBwD36dUERo2c6m4hry
WKgVFOBSSGoFGvrU0M6y6gn2PEWzH6VAgk1r57Q+jHzTVMuJJZmOgiz2giOiJLRH
ZcS28kdKQwZz3r/Hg2/R8Y7qBFVd8mdvzm1zabQ8qbqYM1u2yW8e2y+V2YX1h9je
clLC0YbJ3Op/UlfLFwUBV8ZosS4pQ1xz9yKVQVgrBljYk+2KVA+7qb4M77wsX56J
DpwQVI6u8hAdXKT3es+bWCtON358llbByneTGlV7VLN2vGh/6JoPh+jjYcu8ql8O
gLZg70IyOxddNAsMOlOU2KBuy/Pu6fIz9KL2/rgQXsZVhcJgKfDEgRp7iiQVMxlH
fA2gragibBdqNiwLyzKxXUjfVh1E1RJ2cXDzNOjZkN2ZLMV6etSgd8pD06Wm8G8B
Intlu6ci37sScAY88Fb6DLC0KdpUE/t9nHR2JzILegcJ4EkF/RPaX6zhwBRBFgFn
F/tiwUWBBMXVpj/tDW1vdnE1GKr/3SPK+qPhXWOT70idRtebLxkZgqSGLi/XU1EI
IdfJClZrR7hby7GCoiVgOimHSItM1hG0LXuCajWMQGYXIyUeBBUqZqIZXaB4jLGd
TSdw1sdNNF9oFI5iJ/Wuu+A5tzcIDQv1Th8SSlK1PpGUU22hhjPDPknVm2CnfkST
0DgQVZ0r0oHaeAXmvBSkui38AiPP/XiCDHbpincPxeFQOL60rjnnDu+jtq82eMmf
svU8rXC/LaQwrNeTF59aL/2vahuh2vdgotK1jkgydMjrTzm+PfS3hz8l+OHOAdaB
O0tu6QGMrKVopJN1ESVU5Io+R7ff6eQ5fGjqcl+twAPuKCL5gbzzPfyX5nv6ayh0
N4QZ5Pjc+IC93hbyx51b6at7dsfCz6se2LmdU6ckEe+gysuHIg3JOhbskrNWCDxk
ZacV6AGg5MByYzXsiY+urLZIGNgK81Ap5gS5DG/xUTcG3DO+lcKSSz+sz97MyfNL
EfR2gLFbKzZbUmX/my6tnSX8is1PD1nx6fWg+RjNpLNOOHnKt1nTrepc2eZpfau/
ZdvEwqJEeBb2wzx7fTAc12zigYRzorI4mprengKE2gKcVC1Wf53LAYyy+mWk4RKa
Xd8i+EAFRk0sxkLcpcNdt7CNJtW5mOwGgzzBP2RXAv/JjAu8giy7wSGSs3YbXmI6
vAtmssTz+rKCs6FagezFApXZNRIbxIFWG1KNGXZ0W3HlMjcpAi4y6heZkl/e8BLk
nAnhR1BvXO/TwBK660YO11MEJe450t0FKmaJ7werCJhSUg63yUH+a9bOCpNDz51I
zkG+957fSkEr5DSCGD1AZV8GRmtAof2Cn5w2B0BF2H0BK9PLprhtfrkodXRUXTVf
ZFdTWGpPmWj2TziJqVoRMD1208tWlsM//LZL2DVXTAsXDmBBlxVuz3F4i5MUY/rm
j19DDMHPI3fyTR7QMkDlw/rgncO1IOXuuuEzCZWpQWycfu0dP55A5yr8xuHw2bmc
nrZvVO0nyZFQ306efGdCGJHtM5bysF/aNLoN2PAYa1FE5vrjWbHhVLDBTx9uhiwd
Ubz+fAddEnJ1Pgo8X/3mndiNSLeQ2hl0CXBYqTU3jFQrtRGiOpUaDaQ2OXh1nZrX
scjLe2cAtjSdGnQpqK1TAuEjCDxZcm9MAH9KNOvuwNlaFWUEkmF8v8HkwPti1/q4
rMTpAlZQhmPJwi2sM3sf1I7U3o07KJrt7814ULxC9PfCnsOECp+mU4MqMNUwWsem
HMdMX1kv/R5d5WquLYaFsQW4zpSIzSQmIMqD8+4Ac+oKGiGAXw2Ed+8IHcKPfrGj
l7uRvTilELsAGuVZkPb9oGErPRB1H5Nm288Uw64sBX0awoAp+4eHMPhxIOso/0tv
Aw0FJcZOEWkLCmM5+UeiegyxF02M571Lv03I2lULS0Ib0xG0QjFWCW96uKszaRVM
DlVFHqEHgBR9W2tadXlxyvr6YOzq5FxzeQM8mxnWb6rtkcGp462fDBVmJRJ43f7D
Xs+5KQFtnbgJAmkP30EWoEVLchDJO8TrKGRhtGXDHNTQpD51HG9U3NrCcugPVj/t
UmwgC/19GBXTz0Gr5ruP+wWNLgCZnChaJO0Z/V8MbhSGNvr0CSuEg5qA2UUhrPUl
2/7vSBu96FReLcHeqd/Lvah/6Foe0qvgXyqEz0UopWK80iPw3mnpQyE1zyztqy4I
u4W7cTdt2d0+6HrU+9YW+NjsC2vjWC2fTVDIglsjR7IjVibr+uRSZB/Io5h9YEP4
LTdqXRee7LSyoslG3acg+hBvIUTMonNzCbIjQVr+6Zdjc8RqQbQ6NWkPqsPup88f
qIhjoq2Aq0K3jpifyjcjrMkDeItKfJG4Euum17eK634Rr95M886uoBimom+/p6fl
V57e1tmoSIvAhMHe6Uepkq3uSyL0x+ocKam6Oude/ljHn/IS2dHM2jnUo9A3gJre
sOIX6oSKqGqHpr1TwT0P1o9qQV3R4mlwcPbUh63SmaSmErsbgQuXCLlKEZPnAoZp
V1YuHW/7OFL3S21EhpJSJPf7YhhZSSHC7dfMjW7ImE5trImAkdrVMVFs4GLMzv4F
rv3bOYSOvHXoIBZo4D7NYV7YlEj1D0AI+ygOjaUyJHhNCAfi16HDW4Mtnw/VcAWM
sO7hQuSBPiW3Bf/pvE2YFsmB0bYZPy6KWKW9sIFgMjcL2h7s9uiEv2bPLLNPk2Dk
rV5pVNb1/WuMOiDv8bNuButm32tRNmsHhJr90494A3yR4LAMQ2lXtzoo1LZR/bkZ
84iM12CR/PwD5P50onUtv2M4Zn6SaQfzY+AeX4PMyc79ygqYs+xOW3dtwr77teHR
baPyLIrnVu2ZV3+ZiN+XtVm3E2cZyO1heC426on+0qZHZ5ZvYUn8ybge1nhZASab
+Oz04912grirpl9FN0YKtZzkaLtm2EeyUIxJb2yV2+wPMj26ue6vVj8KlOWRNqUW
mPhHLsicXQoMmwtt7vVMBLf3kq42sj7omEoAHuYFpytP62/4rzeyXZpMxBuLrKuK
P6nZka5PKPMC9yYxLc5adTikq+xHSDaOAOTeK4QSDe2tGbYb1FkTk4TzBiwvnWhu
75JgGrFoffn89asJpo3rK+ZBFkOiEIMLqTBkP0TWhEWMOP7ZTKA6vXr4qIf6aLBR
MNLJCOCBpT9KMvcGEzh1JYsHFv0DHxqY65xTHzA/PyYm6INxox0E4U5pRoOm44OI
sZJ+AybvTRrbm5hkHJAgyWdadAUsLUTsbmIFImPJ3YYtwGs3dDIv0uqR21Tm2m5s
OpYqmxEoULjRAntK0JxygmG/c0Ccbh4baAKlDIEqwhFAsvTW3rqdjl/qz9cQs6Xb
xQgMXGhiUTSaJNHu5r8r73l4yO2UwEx2NE5ZCrvOB1dzqcfDU2McF+2C3ltF1YpP
5YI1DHBVLXeYV4zMp10ueMAqUqe6/js7ySHUhNDeFg77psTpT9UWn+ivypVjPNr6
vEPTtkejfKG4Gm0LrI2Eze8S7C8HgrL2EJfCQld6Fq27ozq/73iaEBgbC+HedIOb
ZRDrdRBG8ERe468NJknSH1asJAnz7veC3O8oNdi2UGrg/oE0AahdE3fYcQN5bHqW
6S9WeBjHNbJQ712LOCoNamEYUKpxEaAYPHJZ3p5v/p4meJ9SXeJfPz93y9jbOui2
9upflF9eh8E6YmbFLOjH6HtrNfZhY0uODqwCMEiT5zwjNog98jQbw32aEMLkoe/u
c/JCR7cyo7JsM7OB0Q9W49tJ9F9j2br5CtRsUs6gd3Bg6GqVgnM9v0bsuYLE2XsI
6xTlwMFPxM2GrMNCrOWppdjtLwccp6fs79MSAZlNhUNd7lOvbR5ffpxBI13a7ycb
WNcpmFZHnQPiptp42G1gNk/y9OEWxmqzCiFY2l5TxtAG4XVw6XjZC+UZfwKZPJFV
hw/icLqxmZ9ccRPbWEaG17uSa/cFwkr+h0AJc6IMSjGuxYYtX5xE0JsDO5jmsehl
z/ulFXAHPwtXIAeBow+WzyOvbuEWrNMCLDtrCEhByQBaMRcjvdxLnrpAo5x2o7Fz
9GeuMTiFMbgHiDUZ+BfZhjjND6PFTtpRvQh1pmJYkvhyvheyfivSgB/Q8g0s0wMQ
6M3oJ62RMrgBG/jiAfdIwnt+3sVwT/tvNVDs1YXFLeIA6wtigrUaF/cdeYttAroZ
O27GeKaTgtp45XStWgRdbKYbfakwDE38IPKs6+wOlaOUew/x961la/lg3Fj86FRx
0ykalyVfGptFOuaVCUu7DxZC+jg7ji1lvVi6XdAl60xHn/Tv4knBiZQ4tBZmP66z
hcoENn/tnkgz4o5UY2iQsqaFltTLKL1gJpyvM2tlChuRm3ogKpO/p/veJzPSwcvd
6fwfwpGGCM6o9LZR9F/QfzMy/YtYwPMR2ysxt7dPT/g8Wjs6FDReikfQZQMA9snB
0K18W2d67P5Sb1V2bo/rQTxlIsbC4M8V1RcosHDn15YSWa/hqzXwtfoU+lahRFDO
QOZb+ll4enHydU/Fu9nkJUcIAhQLihytnQ8ZNrP5yIwnowXKgM6P0HyLjY1mQTwh
FIgOAcHQ61Db+zhJNselqp1jp6ULVmO5W1Zd2xQnsncz73HTtU/gLfY3qM+Wl4mj
qCBC7tkYcU8Yr5J92xLtqO82yWAdFDQAHJXcmM5n55B5fUY2qMbTInRRFzBSd9sY
tjXOyUzN/MU7DEBnBDp0p/wPsf4CUWbgyTjk17MKO2gHLsr7W8kUjxVx84CoRARf
zUMYYAfAY82oFvuTJnPyBNwXnOsSry6cMmHlXQwN0k4BbA37Rm+39y4p9uH+LFZ0
0qCz5JN/rkj4dUTuvjccYH46tpN4GgHcCrU7CYVSeOJZTPtEPnorPnEL1+tch+Dp
t7TDA6JG+05KuhHHbHAtJaLATwk0G9es0Z3LyKvH5xEPoUQ5Y6G96mbgRISp6pvs
O2HRDYsY2rcX4xnL9JrD29CpIEpvRmNyKhGOTq7K4zcJxDNXX/P0ZyvwecY+QIaG
5DHO/3O8CC2CXwrEDkwgkChtkLfzspsll47SjdShSUfEV9jmAcnwhQMOtUgEuO0u
UGKlq5tvG0Sz64klnKZ/orC975UDOdJX0Gw7bKrFJqM2zKYxHIqe+NXmtKLw7NFG
x0wOvq/7noCyDYJ5K3Cck++z0Z1fsRnapmLwi0Y4t75uLGdLbArwWYiRTFZP/xzj
hjJZaWCXIV1kLh5S4nWoPOa45DXzNZDuBJ7yA3S8Rr0vjuYBmxyZa108e1J18Kru
O800kEOkOojp/1v5yNQZ/Z8JLdK4639weDm7kMTE2ju/BLQDM6mhsBVQHnkeDUGS
C8YbIGXtU4rSjXxtVgdu7heBhKmjXedi2oMFeXO9cTclQXjluB0Myh2jkV3D/RYd
wRS1Mc7EGh3NKdNswLRY4LnJjYvw/gzZafUA1dh0gEa99UANGsS/UPhjRkPwjrbu
IGVr5mFOY9PoGFVLV5oiTJVkVIrnRlbmSbFvrU7aqnY4Xua+VcAadGSeSLYjm3g+
QgqRqkulS9veFzhqhHAJVMtV8VFugP5zMQH3FHFA6jH9qzcl/YqEbTwQTEnJsRf2
l0OhmQPbNQ79rxnGRvLfXyf19ZezV16m+viqf+h0A4JMu1tvRFydSe0KcbknjAGD
d5Pu/lG/t32MtxeznBgI6MbIgNEZFSPoXkMkdYvK1dp1x8DJxtnoVKnWf08763a2
eZXwcLUk/3toSKVMtNT2HXAADgvuBJRQGS0jDgLduozzz2y6v++O3kI9SBd8NB+G
2MFNt+7tyUMypoQNLYUfNVCXx9pBmvc+KlbM88KurGS7xF7Xy6+c6Y3haOAxn01G
4hKfgYpUjD98xd3GiGIhO1uDfKa6PFTocFJ9Q9dsXdldBi285cTepKyM/d2Ydz41
Brl5LqBjjBfOmxsQbVlBdXH3svvbSgriLPW13HPJTWdPhVwRrEehjRZW9z82qyt0
/TUpz5aAc/5xaqCBGkqscPLrJJmHPD6aQdVlKYpA5ilS5stq6w7qQI3A5WygCgrc
TM4E+kufRON3ztAc6Vrtothnqrk1550fdA7C3mb5DJ/fNDXonvdyhACh9EJoiYqq
buK5oy3pstLSZPNS/TtgjRB4IkijJJHnEEAiYq/k94EWRMtl3nJ+EbFoJ8XFvqpg
gkRZJlkn93GoCHgls2Nxzw81cB6EKNqY+aKL73NvWIlwT2eL9RmjFzS+sIyo3Swe
FejhDAFD9JBbIQU5ZRhcE95wsdUUjEdJdB3FSbDGn3hLbHb1N1a3XpAzu4cFQFgz
vMD4Y3G10zfk9tNVrouWm29eKRwFCF0VjKbtFzCJcylPwEylMAeCoo+ZM5PxEPtE
ZkKY0c/bt9xfF846Xt5T8RtgVKsTFgZSBM24+G/Mid02V4SpOZblQQA1bUy49ZMG
bTrVOm7nUOT5hsgi+hObf8MV0iFFrIOtyYb4fRSSNo0LiHsdb78I/xrbDSOjXNr1
jkOQ9xb8lB1Ai4QQLvF/1YWvGysO1oSd57A19D1qlVm4nu+q/NEN/zRUGBjGUlZU
sb/MI5aFlxbeXHi1Qie3dIvoGOi4S46IVrIZm4D1vEMNlXDMY2x6/ILEtsfXXPTf
GBtv4AMrUPCAlZCzHG5vowvF605tm6rxoK5N1GnPuq1AA/3Rh7L3oSfRsUIifFiQ
tPZp9olewbupdBZsr6f68Ja+U2dNBOJQMUw0FDqnsQ4f3z9ldY0Cuql0e+z+ZyIy
x9ddaH/hKLHkN51msdvIjYiaFwXljXp2dfSsFOLqajAF6wYGpAtVa96XMpl1d9vb
MbG/A3Cefvl7VZHFpsvMWihFNuOSh79/iOnvDQRucpuw+UeeZcVcorHjG6ujSrK6
fvqRxbRmhETHAsDtU0fMVWZF+IypcZozMZUIHehGJnAUh3sVxFMUC5rMyj/k7/1A
VdnIjFBXcBpxXls3di8s/6PvZscNDncqWHVw00BdLOJYLWVK2EeUZubZyVJrgyh7
7XYkqCgwOEi9E+M+fRiMh0JxN+Y59Ec0uzFOd2x4yqRJryFFuZLIGCxVbE5pzLdj
fORZXtbrZd3FO6w9jRKFwoB+gve0Vc+lW8CHsduyG2LHt1+2Hdi1Q9QekVTBFql6
iFMu1WFfsc3GienwWXb6yOGJqWZCM9h/6zE/Tm03xTS/TJneIwmuCjjPcxRX/Wor
f2HWkT+TJ7CJ8QRnzH642bIh6HIMbiZkPStGBaZdo1iy9XhHeXT36BS7iGzRkO/t
3NIwK+DRhCtUBxQoiKY5RIMSVZK9IyM95BaCX97d7lNWcWibi2q6d+RIa/xQP+Oj
kfAgAx8+hFlwgfwRb+lKpf0MpKfjONoL3sGHH/sG0V5tJQF03ec3Fz8N7OdwWnRu
JXZaadWpeDx0jXeCyo81WlClfkNaforbNHcxfj6M+6CmpLeLKnREN+zbzcZwb/oP
tZSR3ZsU9L3jwMmcta0lzukam5mxl8kSSGoOk4ockakNx+JtEC+g86n65/VCbdZN
mK22Lxe3BlvfBMdmzVN1/6rwZGjqET+1mjOinIiafJN211DFxi6Zmye5vHL+nzvo
nLYh/Ks3pSXJAs6LutFOOOUJ1bRcfqkVeZUseqv7lY0asura+Y36A7Uas8npOUvY
X3UBGc2dXRKjMnAUUKEPhRC0yvlPmy5TWKjOFEYyuy/oEwJ8GC/ZL/UWGGC40Ey1
fHToJXo5KR1E4dPtBcck4CZPSasYvOxuNeZlI6VvuZN+bS+BKkxo8uc/GWe/V+k6
5zoNFA6u9wuhlxQ51G3YlFahX4f27HTFTaxZnpY/dkZaH4TM3Lo3NXvvEAFJVawX
aJwE3PDIm8BjFMbiixfh2ZffHUt3pGCEG64DdOG31TYy1Kgrto/HCj4QqvIRJHUM
kHU704DhJEDe9N4OnHZuNQbJkwcxfEXHdwlzb5moTiIyS3ETtUffX99YxwnzVvCi
FeUHDSOb8nOUHgX+mWziAFAmFG2wR8hKk7pprpjwMH1Mr4L66WSIdXCeqbsMFEvM
HowzwG8/4Fd5uRnS+3XC7DmvWC8/nb27/hQ7Ewxtdvt4faiOzT3wXgzTXU5CDsPt
37uEADz/rTWeOsKpRCupZpT/Bks9BdlxQpZ7hjpUf/uk0IP4bkFl8k5+IvTDpuly
rE2Ybxyzb2W+aPXLq7rSR9l+vz7WWMc8NYbA5VleYojQNoXEMTREoAVnIje01rOa
7zWt6sEJQIOROBi8fzwH/oQWCAtMr2WxOj0p4Ra5DYCu1+1SJFV28jpwwvabOcN1
zFkLf12AuiQlpdOyxTMAkVK8rrr89a1mnFi8o5JqbavSquIicFBZupkYXeAQReNV
oVEqnatUXMaruP4UAseZCaB2DOqgeuAdbKBawm2A+kuFGBWHtiDZcL4ButnarGGw
/VlXsR6DI2Q/cf/rN50mCj+h8V9g1gEMKM09GooJA+OojDIWd8V5XjEg/xEquG93
c8OWRehv8Til7DYMZa4r7T8TlaIaRGa6TOMyH6/d0KmuaV6NJxr2+aBxJ1pIThYQ
4Or8xuXIM9CItUwQdS8IkYF1QQqdjasc01mhndpolaRvAigN1E3teEFpNdUOfDE9
0ycC7US2PJQpKdIbMAvNNDY1x/TRC3P2ueVNK9bZDYJnGwrpsUpfwBD0R1r4eBIZ
Gk81kvEQO/8O0zx7dj0p3fDEEQ2KorNJTttFOZZVqNqTurruSHCY37GDCZ3AGY4M
D/jFTR10z3Pt+/y6M/zmJPluXeK9BZwlmgs+tGq2lOSIzIXfeZR817LLzcB7LBBV
N7YQViCeNdMqqVG/a+hjmfGwFfZ7xVSgy5qlQLtIZSfZAvtl/9CmER1xwxFNIq1U
gKjVKaFzM7OpUoieF0nDNARvrPV4AD384C1r7jNebAXKHye9FQET3+d3dD0+D+GD
jComQwhbV+Frq8YP9PNBf4Hp72kYk87J/6njWf69gS8BDhFt0Gu3jVrFzQb6O7ur
Z+zGclmQF++GG2nVW7jZohh5foUh+ZNXj12G6CCvf7TY8V/41+XUiPDAxgRzLHl4
CgK+vE1kO0LFFoLX0t41fNLOR14ipA6G23QPQ+yQFtC1mlw3c587akbE/i52Izw8
B7vweKPMIUeaf2eyHdebBX103QTDtDAZbKeXB2hWNQSP0a5bOAAZhEIDHZabX8NA
0OPHH8iKZ6PpqIqz9NtsvG7Xx34RfKX+Lkl9+VzxZz1wOFY6LgP5ioJGVDWWE8iF
RHMaQxeRVa3+Bt9h4crqPAVefSyRcYvtV5q4G1hH48OWdicYslkx/FtnN1hwkkQE
IO6ZT9T2KA8+dV8S89mPYn+6I9zDi9t/7hlqPMiHNhtD9QLZo2pNFlkFW6c5HIDT
zFSgEO6sP04yEPlaOhwTUwY9CzoWF9JE1Ot2O0gEp8kSxpvk4yo9ty8RG1V5/qIh
CrlaWsrMbYg4qurCUDA9SR3iqX15LjDsAgSpKh7F+ScE9v3av4V3GZ9fWRrl37lU
5+AQ9b8Py5NV4Nqf9QHSnTGelGCeUgrUVISXSiwzT1sqQCloG43iK4IYNbpjnqFx
QNBMfX7aOfuZ9K8H8D62Vi474GHtzxKsTzjNAiWlO/AzeNKpCsLZ7hgCfybLnWje
zsURuiVPT6dcxIhNqudyq8oZf/iNmjBCxfDanyQlvw7NzFlVilXptkhqo85CS8DN
Egn4tbIosP29CLZgaZXifrmHFj96oTOPg9w0d7z1HlTqfJvNyq3TO07YlGotiLqR
DL6qbx/y1DEWeBNvaCAx7cxtMyZ143LxDpGeI+de2aulVeiaCNCEAaQ61NfuJPTL
dcxHrWBlB1BSDD42QJX25b7F7rkWDqpaumBU0gJClnBQOvhMfJQFteZz0ktRSwzJ
wgIZaFKutdZ/9b9J6ajYrwZG/uOAyn+A4U4YT9tMK5CYJxAnQXx2ykzAAMP0xNJv
4uCMyRmDZ6h0x1ZBPtaaU9OXU67SH1Hpa/mzouXjLUHUcHNSwjNpTYMJjXEK6m+m
MS8BvxvFjISp7KriKC7xY3r6XtCSwKGnbQyKjiJtux3SNg7GOrQi8Dk2rx9z9moL
jFIguBzwBwNGV/ymI62Yap4UWBGEcl2zXG57Va9gxlfLpeOrNwnMeQ5Mz3NcbfTZ
Owt8Xqhokrdz6WYFYWs0GI0hQTHRtsHxaWu1v17BMTUH81knYQ16jrn6tyJwB0Cq
kxp13LThmZ5Qsbd5engcfxjePyOtp4AYrQfZIJh2cofvCZ4VNtWV870/z/ZditRA
7Jz8TiZrm/4W8tj3PTfrbho0Mg93r3VP8U5cLrMFOjxr3ynAr0x1SjI5S/s2FhcR
lqTC1CXf+h8QzTwITXUmSbj6dDjMWvnsdkTHKxX8pXG71NHyylXEAGg5OgCjSvEa
D8EQMWXPCxSC193BrrApkDQdtGrXTsX5vfm3p4UH5dKy75rys3gCjO3telJZoim5
IxBBPhj+2dVbZ19y/PWIF/7LOdeI117KHXSq1Dup5Fb2FbOsfR7N/0CP7VIY1SJr
FVwdNhYO04QM8neL8Ikx4SXIPV+UWK00t9zfVgv3OnnDfrnOmI7CHBlLD2Tyuy04
qy4O5IoFIayI5YtD5fpVRTF/7JeG+XHupBh4PH3k0CX24anANPIrKGFHCp8dfDv5
J9jOJ5tlfaPUpCJBiXFigqUrf7TNzVDcl72toPeZxDnJGjInT8xjRsX2ZAm2TGVn
E+CNe+Ve5j3lwkCPN3/2ela0OjCZ731/bKtcZN3u8hj4oxzR01JR/8TFsWS8lRlI
DWkTL/uACtP41cJ1lkcVUyq6JYKrnbjxfHC/2sdpKg8ucs6FhIrOPGXxIZCmjDmU
V1e2TYjWJthKx89RLZ82Z1cu5uPeFuE5zI1NatEWcWduXp42eyC9UtynUEtzglbS
waGNzzOUjZjnh7AUk1P6q2NCA2KVGJ6TMGU39kBIesSoxN51IrQWmayLDjNJz+qH
EQRRk8JOMIV2rfz/mu+BKf5rMrinGFFa6bIMfyuFxWoGJ5lZ4nVsRcf4U6rzhbhr
iQBZ8tVRZS5ICjFww+HMCoD9B5X/pAYHIhyh5C347owW4t1nc4iUCQ4Riyn2JOuA
GMHHTcO3aoXCCokMw+ptP2tgaj2jHO5Mgjwid3wXhumqgzHsQuPRiBR0kRqTuHvJ
w7I4JycGZkuITyBu2JrgiC4kX0HcauThf2++La2zg7NIpI4FIPRi6WzbLunZsBC+
nY1H/bG9CgVXCgX8nORm1zxqQ6EYY0itjDM1aQgqpeVoTZZQ//YpHThtZTVEL9Ql
ABygmspLUUeZzepjN/qZDqhZFHaL19sX/t2UzR65ameuhvlreh+cBZjnFwe2ZPlt
WQjcs33rC2U1NCE4xlkR5b5w7Um8FPv4L1Mi/twK3moetqhEAuJxwuaXtAFUPyoC
1Gm/RZnQyiz4Yxhg/FRjaWH24F3bQDWc/LTtaO/xfzgl+0OabNiOg7Y+FUOo5l+F
yRslze183Hk3LCnEMYvhOmDBNPv8mcfriWZIN2hovsMTMN5RH1Xw7hEvDvfh127z
Si+1pd7cXUBD0cq1m3FZdADJzm5YXVYwkVtIYvjgFsHei95CKUxOwePij0jkObSh
CWsM2GZlST7fONEPGbAcQw3IP0lpGVsRgTSwifpa1fZ6RosCFgmHt8jolyeOBOpJ
7Z+QFyqw8T7LM52u1O/6ifiltj1A8+p3yA89D9HbB1itHuIHScYi6awfycEsN/5z
3AQZW3vV+z4oOuGJ6Dwv5mDys240EgiyiESPjNT0CU3QtUrrPrQVrwKVbRg6sRV9
JCF8mkpJoYWtsbvNSjVg2WbAtbBi3DtjSmr+5T+aUydQ6tapJ7gM5k828KUhvYC/
P5h3G4GLEN4lVIKvQibAtVUVuycRiAtsR1vNsxGr8uE4qxrr7jgylJzTczc8TTtI
L0ZN4+KQcjy9ZVXwoJ+5tQWHt3GWiihVpg3SAKW+Pw+Now3Cve9Q4whtygFmI2CM
KMorIonunH9mcpG54fYMB9wYCkKNpsbwzBYCTZYUSBEJoTc/O0JXxMVc7/K/XXK0
FI7/4n29lYAHxB+166a/2kQ3myCoQfobH8jgfuFfjCFNXuSvzS7IF4pGl37odhGH
tDkSOejX5AqtCoUiRxFLf9GNqy+v6H1rr43MBchRvZrMhWY0WwF6t92iicsoallP
vAr319HIj4oTepWp9XkX5fHDydxXcA8P6OeO3TACMBnd+AJ6A/Y31TYJO9T72Tg1
5XDLos35PGz8bhbVbMc0Ra3Txt7knrrEdkKeA9xyF9/BKQsv2LKoHUHDWIhwrm7P
xcrSOmUdKinbJjqvVaHr8V4Qalz3aWtnjyLpJT7z/d/P2FCQJJNEGWb614Lm8Cfc
zv87jXXEDkL1lWCIOUTTM3M43TBAy51DGSdN621cxi7UDgZP1PcfyS4cplUbfVqT
HMDsu8afebbJh3wyiVZbdibxs7Zv0VrWZmf17TI5G4YWCcbmq/lGYTIyeV2Joj7c
DT3KDX8huYkmbjCTX99Jynu6eLEoY0JdAoP8GRuYAldwGpZ0JhLavQEINjn4b91v
A1O/URKkY0ZDOoyUPO8UlY33rsq9iAbNQBe0b4uPeEzn+Qx4APyLmgcDw7gHKA43
Nmgk9y89cqh+KsxnnQjYTE4HU8uoefSBY3w9L49kG8MtyQFYEisi/qnEUl1/AyxX
uAFPhGqjQznCB2DFyBtDKAj24jKSDPT43IW+fgR85ab7mUNm8JcByFKfGDVji5Mw
AWpS3UJ3JlvlglHqK6er2FDU/F/5p/RGIprZCiPpOlLQpmsL3cBpzxlf8h40VVyN
WOfwHyCaPoXbBmo9hEBDJW7lAJE1o+rvCyE5CW/wh60/+w5purj7Q/aPmVxXCHfo
9PYZOkBFAbd9aNMx5QyBYk/Nk+C8FgyyZf5jLN5PxEvFU71ENAYnOCRIPZAR0UN/
GxtvGHz0/8l1RaI8BUb8DcFB51fPArYwweMYSZmAywRsPb/V+9nP47zVljKR/9xC
zzK2Cm/+bnmwkEHVnQAIyqE2bdgFGumnIK1bKddl7fHpnn/EizeAmAG5TtFChK5c
Po6FY3L7GSw+rfEemLyqCmA3DtcIgfKJw4LfDOSZErlxAe3AXpASoQgqQjVJOW5J
pmT6q726S+n3l7nFPBST/ifTK8kKarmtCGrcpPA+cXq5ibUTKVPVV+qj+iy1D6CN
gcXO0e0A3xN2JruRYbjISJBso2RRntWRzWkxakaRgLKovAzixP5yP5l/2O9KaHaU
dZ7XeDtceW+oPD5AEHRSd3cfE0zd4UCZdJp7aXpnKLkRvzjnxIbD51tmDqmYdVxS
A7uPz6Max5OzyN0Jkk65oft5QrhM3SmClB/eGjK3DXcZLvsQ724U6D/ZiBCXG+TK
OtRSsilz2b92APcNi/lL8WxDaQWY/lw5T7gIvIIteM/KCSha2nljGsGHd3smE1Zo
Blycu8kgMaeyJZ/IFWIz0NuM3bXVyxthj9R1fqC3ZjNCWPNAeNYh2ZNpn5JMLW5y
e6MkpIHzPLecQ9ScR2Zj+wo/F+icbMKIULE3aOEFz0xxEe4Ull/fAxplZ8s6B4e9
Y44gYtQD5pPXgARgdkFUInLY7LN1SQzfFmR+xHyMMzFQX8tapTyF3T85Du3EP8ZK
sbIpLTvm/PTjp7Gl3f4FBICqglHl+yamAqz84uZBJSHNonUiV4woAY4QX3eypTYt
VRHXQ1X3z9tdj4kQfmCS1RiumU0hriILTZuGHc/wMTP5MK3EBYTuWHh5pUCymtRu
tE0HzKjO+cuVAa5KYjNEYDvyCgq/pXKlt0RsT/rBgA4cB0Wketyu/0PU2dF2nEGs
P++JOxNsAWn5e+C1sJTbUogWDF4agi+IaUxvIS5S+nqkqMMkbvLpYD+rFQeNyDwO
7TkU1Gg/9DQGLW6ZRqKnhmMaUTsLAYLwo4ZOqx7xhiatylN+4KhbVB9n+WC+x8U5
w4CYPBNjd4eu0Le6T3af4px7xhH7NBvyh7maRNMiFHqOXUqoUPcTRmGA6Dgsa4Hi
o4WkuUi4L/Uw/rYMOMkDsPuzQ9o+jZtQTwISYK0gFYqqWS6zDF945ngzTqvIYsr+
mm+tsZiccvMLMo3bukNIMoKSSjB5ZnH5pcZDu41hyiMsLk3BkuEhi7UZMcGe1znX
e+Jgd1H5G5/BA24Z2O665yR2zBA7QeMmAf/7z4/7S54+Y84L9V5Jnn4s1KmUrsmk
7+GE0i6WtHFBPjCp8nNy0fZ9JGgB+rtXZJgnRQN4PhbSwPKaZk7GyalABVJZjX4G
aHBSz5AZC7KoBjABCgSBmlGU1eZM1HZE7dOun/5goMQy5s8vxiHIpl8jX44QIdmF
Po55xAcfj7gY0jNgHXOIHu76fL2rwH8F07ND7HepnVX/QCgbYnvL9lh0HLs2ggSj
2nsMMVSAgQ3Jzp4l8blyP41h7i61lxBaiIU9ty5FsWABVQnjDh38qgbbJHIBW1io
XGpIL2/wteF1tq9N3UlUjGaL2JSXzFsxeyMnFvTx7ovojXR1LCWKDBW9u2VV1/uo
/+GueUzW10esAIAJvd4zeXKISTBlqX68BV95pLnv7aTorNmgApqUHOzREersQPD8
Ef+G/drD78pg6ICCd6fPhl5ILdLtUn2h3vWZKtWgkowR7HTgxKjWPyo7iKTsXzfA
8SPEqaS5Ny8VCT09C+fjXOnggmRN5h3NU5ho9rfoF2SavCQqQlSRK4rElQaGbmk/
2p5zE7CrH5tg3AGHW6X2mEjSALCIK/81OhWpfjNQ9+Gv9V25bZj/h6MRIZMit0V/
F9iCVInZ0XgfKSjHDQivjA0lkc8N2BhN4WN2Y/goIz+943tgKX05Z7f9rcHjmC8M
+QWU8hbit7sNKyyiykjL0Kx9CJAQN0M7/R+1HpcxVl6wGwYu+hwdVs3tFEkLUxBO
VUN3aYxhJeMj2q5gXk1ZCKW9dTHHvDS4z3OhCvOqDonRu2htIeWCVi4QGnVb+7cy
MxVPimaOUYIr7TA+MXnnO0kEZOE0QHS3fS8gMysNULRAfIzg43UyZXZ6pWLXnxjm
1RDT3Xv7oAptmE8byHORSp/ZFWoMo6Fp8s0gur1d4QdxbjyFS6y3ZHXgmS86i77C
q4zg4o5MDUwXPghWF1cGE4FU6x3239U+OkcbJje4CwsDShCwDTFpO0zQmH49kbgb
JH64CJh6yMHGbOmzGbfoXMupynP/SyCLJuZyhEkpirJV1DO3i5HtpCYrf8FTtw2a
/0DnEy076dn8b8gNJXF+f9E0jQkLnfPe594B8P2sP6SeRNWx83f70QGHZtomnGYL
87ay75FpQrz1i/F6yX9iLz/mjzSOnF6JXyxk84F9xIw+ENq7dw7TvWmNkxxaoLvm
buvahBuz9gwXTNBwtOjGj5cUGfM+nR5zbnZOr+S/0A61QA1le6chFK3+JLwYJ9oM
9JvLajS56Jza5Rt265W3y6/moZZID+ouIngBlnZlRibfcGLHSuvhbg2IYWXqFgid
UafrrFNSRToho8WnHfioyBFCnMbvIbq1ZlnxgBgCKllm0DxuZKlU2bTUT74Rs4EJ
v9nmdDiyW4/oDnxv8P3I+Azpl+3RVowU2f7fYez1NHhSE9iuSTVt3TN2y4EsYVSP
Lb9Yriev2xfRGOQKXJQCGZ/+jcuqlfoFPrbwRDYlUFfcPrW7F+eP2yeayY882o5K
0o1FceWfHKwWif3cq6eCC+mphatbvTJ5hHZFyODuhPnYrNI1GjWVLyIrvNUIRGRx
YclpRYVrvFYjCLoF+Jlujj8GrquQmIsrERmSPcp36LMeTMmaN6bjDktJI38qRb7U
eCFIsBhD3eEvabUE+Oe91NvV81Xepl0CrwAA6Ot+PY68KK4Lwelf4QX6BbbpioQI
2klsrrnyhWq0yi1YS1aeajbJLmloYVBn+yqbP5TKB5mx4hwiLD/xYg6bxB3wE6GR
c035gH4mWsI5Xkrg2/v53DAVstLNhxQFSn6Xk9ZqKDOqL/GfY01/vZC3e7XunaJj
s4PyB9ppiTSV0CnF88gYrLTeCYK1msEhlqYsvrOBt+UzhL5ETea6qvO4HVEniPY4
qzTeRgPphwdUEy3UHTTl5TdIwRAuCsSb56M/1ObVjxhwm3sQPZDscIB/7pBzLup7
bqrjjmNAIrgTn2NGrbGR8CKJK0RfURmZ0qn99wa3Vhb5Vqf74z+Un+IAwoeKMKqW
AJ0xgOlcqnJZH2fF5VpNg6ljpyVhj+l3ygynyMlrZQAVM3oICfwytkAHw41JddNd
bbqCOVyq5W9s68pgN7r3MNxbphYRGM94kEJZ3/3wI66UErQbgcpivBafn53807yr
x1IXbAk8N7JbX82s3az6h5GagAHSS9bYEKqFlwJGhlw9HJ3+Xblox7QnfcPKqjIT
A25AGyye9nmSQZ6N1Z9Ut30d7uLdQNngmRzwdUQj6s9l/4QuKJWEwxbIfKYOTIWq
5cg0Yt46e3v6qwCqSslOdK0ac0WwgEDcN7aHrbsiPYjopcGRE5sIma/FEy5AazTh
bV5yjuqVYmnzxY4yeNWm4vNgyTyrw2rBevYYN7L1eCGsYU/kPoDfsaXzYQIUhVkW
1NVntWmrvxrjH2LPazEQPGYnJIHtPhOMGfWQ+dOBuQejGHbKzAQtMnVFbKpHRRWy
xLbGo85xiR/IFbQMg0ChtHFPDRmMLFVCvsVDEjsu1k+cQw3VxOHOIVnXlpMD6G3c
SyN1zJijgdf0Dim1E+khs6Gt0dd1t48pN+eJLO36P09ZuuPi9yRn+J+GzjUn5XDv
uphadUHueOS45JBVTaHCUltnCO3WsY2i/zS01StJ1ee06BVeO76Qjp2qrmUGXU97
wVbxf4WlmnmIkTjkvdQiQB9A/wB9m9FEbXaPHm3gwonTLmuIm2WvHuXeJRQmB0l0
jl3H9zey2GjWRm2AIqauWkAphwu4p6RbivWQ7seUEr6ALvO52UuD9Zrl0R2ygcIH
vndV6nZjM3C7c+QP3ArKd5oguS+URIypw70Bzab5lfpOz8Zz0kABU0IpHSdD8gQA
Lhg9AAYosq57lnCTuno20QPB+zmuxQyQzV7+xJIEDuOQ+rtJDM6riR5L3Vgzp5cV
YmWRtRzuhUzCgh7pbBDMNaK1Ee9TtH39j8RiTCbLuU0edFfX36yCDGJ9WNfbmYKH
HWIOyZYgNX5XC/Z/CA9v+JHdiF9+MrwUdQ/HUfhfc2nNgoDdfyqU1zKtmDQ1K3v9
29ohBhEEq8dKVNo8XCbSZJ80l9wHY0KwqAMh2zVMlxFPtDTeTd42yT9Z29bD8oxp
EG1Glrteisj7QXEu+MnAswlbDN8xOatuFhuNvELT7g5nchLzy9+do5Abp/QFFz5U
nFCx8RG0xyJIhR+8n3ezdYxD7q9KtccAY3ANFFVFE/9+8vKIeWdeCXzeQ02UeU7W
J4V0sFZpenc56O8Jo8tZgRp3IO+ZhS02/WiXwWLL2Wvl9h/EXqSaUqn7wcGRv9NQ
gz6nBYJKlutd9OSMkAx2KC9yq9AT+mEmem4VeU96eq/ffLZVVfRIJ4JIXuauiS+Q
GZs5wewO3Uv86Gw+jgMTXufYTFXfuQ5RaD0RWTDGSh0YJi5R3ZgsjG8AEIubV9Td
1p66n75zDoIQaAUll2t8N3my5gcKEhwoOlSWzTLdMosUnjWQ0EZQs76qJiwTRTgk
hV68U4Iy5qIz6vawmerkGUFdF3QntMk71SIaT4q5bCOUhpN09OZ8BXu6U/U1bzKB
//9nzFYwovzuXWBHYuUU0fvp7na/GYAXF3CLoJ7GzpmNnM9glJprRydtcw3ffNkX
ODSfuOIhe1/ncYq+Vne5I67yEDi8OTQABHZgqSmBBSDwwS/OdHJeSx8LSOxGnyF/
ZjcIJGKH/IJuVmOUT3DOYAsjrkKPu8TlQbGn0puR1vQJkGMYPu5PFfSLPKNpFA1k
8QRj9T/r8aTcLUw1UgGTAfPF/NywwtKx0nV6+lQKTaAY6tbJrJF8f+Ot1v891aCR
gTfBSHsdJrT7wdPGSumqLIL+BjDx85+8zKJbd+HJqtJ8y/DMgQ2bY4Qbufs1TH0d
B7fTEGnfJE3O8v3b3sD5NLm0hYZP5sZeAW5YZYg1S9ERznYwbP3vIXCkFTCFiIUn
u9d2MTiVe7kXodvJae7RusgdGLiUqqPKUc2ZW5iUwcz6jCx/vDfXne0xw4ajV/oU
M1PSYpUHw6z2DVUnNyT+uoEX9MkEyjcFgO1AKEdx/YOjqm9bwyuTvOTL3djda4dm
t5ABtp0FrkDSNiEJ6ulTKLd8MGhKIyXARPAMSugndyfXLt9fmfzborM+txR5Xf3i
4SAtN4NnSR3zXRCrLGeue2Uz6cKGhaHauo5Hg2ephPX4vkh24WDNLQVJbKkrQdOO
8d9JMWTDvs9AfkoGGmPDFaW9hJg+BBA2CdxN+Qoji1Al0k0QjzwIXLipYVrVY9gc
+GKB8qJFiI7TSpwYYJNcZ6CfsRNWzG/Pk/Yd4M6KiKJYHXUOIxDd4fYJ7XcvQrt4
6sOq+EkghQUZExPIe6nYXJ/1JbQA4qYH6JZWcv6vNFsqNvq13fW8YB6HU0OInoOz
xw2IUkZ91vBsdIx/Es6QIJZgHQ9Swg3n/sqKalYlKg5C/F29cpmYzfN6PY+Xr5Se
2FeB77e5Tfh3xo31nINk8AzGTvP2uz97W42oPYPeKuipTzYVoByKyeAYcSZIX0k0
SieCB35VJtgZuKoY/fFGtUUN8jSlroYf4LpQAIhf6qijc09cK6usmjzpw25WydyF
OVleSI0XMUp3XK0wcxXIoPnxp6TrE5vBrQVuRcHoumJ4Ppzd0jfupxXeCVqjxbl1
TAn1+L3fGzZ0QIN28XerlY2Rb1WuAg/SUKOcQRJ0/U0xcyGkquN/tItzt72pecb+
URIdi+RisQ8K48C+3SV2SDg/t6VwxlNi6Sky7ISo2SNGoPr3hD0ZeNWc2gHAFQkf
rdL5XfgeEs81TDI0UHHlxSima6kLkq0KpNcTj6YARjq+yYiw0F/KXzt7ycXiBdNm
EYYXFge6/7XiWP/O+LOwINyGsaiGmInq6qzMpRF3bGt7IYXG/8W0Sz6xlr4pICNO
F/UaoY73Kr4HgthVx1ORasrSpw5md0+suF9Jmvsr5qmfOdQto3fgwV2RGgjEG8qQ
d2/WACuxjGOj6Cy3qPol6iUWpxNJj5FncSV6gWW/GbZsB91m/8MR85n51/3UN0jE
WkHnDo4z1lBgNtx7Vsj9zbXVJkuXKu4vj3m98U607OEfVRMOTZsCjt/5xKIFEG8W
+Pma6AsQd5MFKY/tfH7drT1a89RfhY4iCzeAqNVACzGdAuXEPd6V7VU+UrNwVee8
X5CMxTXVAei/LE/p1U9FGfo+dk+MK1i3FkHYyhBpFmB6h4o6wpL/7T4innqHS4N3
SiIbj5FTIBphqyZFB5fMFdeTs6v38/LTjqqTLqoFvhcdtiq1QbDbqD8H1+txANAF
FmIWVg2Mo0Bj3UBKiyhTY86r7nKz8K7/4md1VVF46UzH73eayvuvPFO935y5vlTL
7u+DUwx1zGOjkXo7oOsVaOG11jq/s15ucDovS6sBXK87txjF6kd8cE2SjVwtw56u
yv6poJG0QFhUz76nPLiLmrrHOTFlyG+gpga/tykX2DRlVm8I708yt1KZjy+r6yBc
9hoqDxIdthpLeZhub9XJxK5s2+HhCxUGjete1mZSwVVJjbhYSJPhdUWNPiLEBu3o
KMw03xuBwQe0T7WJkPcyofWiHAG81Fg/OYkdJmqYfVz2IhX0tDtB3g1Ika41rSfA
jF6KbzflHLe+IvanlotiSjg9eJps+RavYUYfGcn6v6hp/rfC6s7LdXvTlqYzyapU
k8ZBhl7fI8PeUsWtVQAec+a0A3xSUekckei+Y9vyOrh1lrmcPDrTGbVpjDs78CR3
/h5XEYENSMKpRh0A7QIXpqDfB6sO8zus7G3g0+1l39gNCqkJeJCeUiB648/xotlk
n1+bdn/9eejMl7AulqV2cGWk7HT4Z2/YlmZASivuVEpFlmNVMOljWHhRMdhupkw6
IbmVd9WZXhLPH/qybmBFfnUY8UW6yHDkLjF6yrbaTP4WijskgJ/Osq2zsLUGMY11
voqS7BhHU+TdwH8Ozaw5S56cJb4HWWI5k/iyRErMq7kbBOx82wu1QZIOiSPRqv9D
i9eAAH/PKoQMgNC4rK03HSo2f5n4sbpgEx4hPLWQCikfQ4WVfEWrTNFQwsKBTzXp
/JtM7R1mH9x/30izNXuxfVDpImuCrnmEm8OHZcJq2vtlA7d8wG9QiAIexXWW2TKV
sNi52kY3iJP1KnqkHRwd1bczmaU130rLtHHJ4t0nKBhbegLKBX2ki75j62YQcKkG
5Lb0GSF+xz+DhDCEJzrFdjK74BPga0XtMsHHZWzNLQnMnE+2qNlxeHaS4hL8C4Pk
cV/XfmklzRkKiGWzWDNIZ7PVzjWCxkVDgINeKdQiXuLU2Eu0Evl4MFzJYPXWKW8Z
3rIzsQcC0sJeMQ1FQANoWXw14EeIN5L/im9Mz5CunTdSWrg7tedFGRmJrHzq3A7c
uyPY2pRPvAknY33kEnw7lT7WLyNHq4o0g8NtZPMrOaXr99x4CjRy46OeIw52uERZ
w5xMilfjT9TZ0TPDENhvt9sodqaUfLQrBmL0F0O7FmxMEFRYban0I97sF29dp7/a
tTty4OUCbaX94VpqmBx48GXUlAHqHHCvR65RgRPdV5VVU7ShuLxFWKlsjfh4Xu0+
QInX1+jbaqncc68OWTjwJrhCvrV0ch4U/oc3JNYktK9RFJBa/alxkA9VqG4Zie6l
DUFLX2hA5w9qFz9H9wgpgcf0sdI1vIeRIWDKmaROfNJk6PnE2aNRq+KeQNS6inSl
UAVP1zJfdyy9hvISAm6CNdCQkyKGT6hQflcjAnmCrfmklkZqagIbT2cGobz9RhNL
KPeWskZEuhgEch6vXPaiIhKqLBbLdaLDftAOMvAy+uOWdj+2fExGyDbNddmXon2l
BkccngkdtgdLmetF7+l6J/ow/cSJN/GuLCHZAlwcU1pv1gzX43zWqXx/EPTxV6Ir
ZO900ouQFyBnaUYfWpNaqMQ6RYC5hSCRl37ajbtVC/XyLAk0t4IyhalQD6YMKvEc
KbmaiqHt1rAU5NYx5XbM5w3uCJrZqqe4Hipg6D4yUy6cDLjkFNcYkg5E7L0idHQo
P3c6L6ssda2m5BzAtT7NKzSDQyd7N64b5LqdtOklJLhjIB/qT4hE97MCrFKS//X2
uMuU1t6MV+iIxM0CiYAAZs5BoHFLLgEYLa5c5RWsJb9TTbIPfBlnt4zrbH24XOQr
E9o04rd3BZh/D4wcN8SfS6f9gzNI9udcp95+IoDZtI9f9GAneJ8VrHyxn2TXwphL
PWH4rYMwWzFqtN7n5OH07s0hHqk3uZrKBoR8ZseGEk2s0ygqd8Au31OIfA3j9uZ/
QmsWzG9nxcOHxjzWOaTmbgKHO7wCUdUsLWaO9uUFgLRCffIioaZEU7Kpj8UfYCkR
7KC1hq5PUHiWW2OTZ6m1JrwUvmiM06byuSXXJQEbuulBLdrimKGWRszWqoq+KG3m
DaFRTjIX0h75dnJAXPsyNI1SZg9MbYY868bEEhv1OA/fu3uEIMtic6Xqfx5ARd04
qhul5d6tvcrjaMknDMNIFRlaxIjwKoVaVX+zkjttOegTlMUuVmcuvH13WgCHln/b
z6JXkL5wwaS4RJCVGMIMx/9O+NVPC8YTeL+1khCykUG14KwNSzmPkkHJKGq67hnY
D8I9QcNuOV7dVZDaE9hADPElSpuTg2RGpuiB59QQmmclT91bj+Ss/7XoZgmIdChY
mwVotouRZ/qtqdnc6slnCjdrFV6vl0VNAO8MIqRNyn6SpyIt2DQvCabiOtI+TRIM
AuNhYKnLxlY84v6MquqhShjQVbpTV/J84/cUR/OAPOe9KsE3MB7GZ7VDjHjm5ZSx
+J3sAgoQC+quPiln/Fd+4m1i0hQWVWPpnWiPsE1tL/H+cejNYdlNFxEyDlYmglZM
GZ6RYPqqXTq1A+xjRbXcjzX8XSBItYmk6uzdKc1Js6WVobNjdY2Ik11b116PM9o7
sx5ZMbL0kle3g/D2CheTysMWTydWmgy7JQM80Z7g2psWHu8D/wdTWNzlKMApfBpp
cn1+vQFuPs1bGISr89uzM3cLLlbiQtIW0XqkAlqkDhOv6Hy8ECf+pLRhIKINQI1F
AkZ/v8WRy9flG9IwVxlqlvwpPJqsuN1n4jQ9sBhr9ubGdM5kKL92MPMDOS7+Okq/
vsVdCnZN9KgSRgdjSHUD2lTaa2Iti6tjFgpFoU0kQDEG1eqhGOJlOLEa+x/WdGLx
P7XJvo9Ip7D1lQBJEsXsE7SejdXGFsw8BvhWwColvL74MLPphBYPFJ0SDoMhwWWG
2aD042Gh2gIp/yc0+JDDi5q5OszQtHxvTyTxQdgONmE3qPIK5J9ffJKsG/+yQ7BK
qWHfRMXBxRM35evDfjfaITo9y25S6FRKea+TxVZQ9fHf9dzOMapNr5RAm2TavIZK
k6rnPV1f4cYXmqBanfiisQgiO8m769aA+QifXSKAO70nN9CxcoJBMQMA+4/Yu1V9
UAGKnhU4zab144i6fCzL2Sy3EFbnhNRzM4bq7D4ivjq3nCE39py/kX5B/3c1jseb
sAOPJZGrNubZUaHrV0GTGaYQ61fMbv00Q4j1Nl/lmClOyLsOS2mVbbddhKuFqkWC
6UERE1EZdYnGvg49EZk4OhTt7iWfqKbbBmlwkENfFS8YFVJCJTg5gkJLgVvtdodK
BCvwABsoiFxwJVBmsEV3muwAinj0VmB927ZKpaJGmA/H2uh6u6qqS0/R6qAUXOjl
UqSZjGZHzP8VLOnhyLBNSgrO2GGHgyCIQUyzT5jE/080wXchXeS7M2FDcaciYStr
x+0q1FEa1Abr2TGvLllZOZcqy18lXE3MAcVwb9CPxm9G70WFshOT8FMrG+h3Zq+z
Yq/F1m6mZYi+No59Kf/cSpX5aHf1Z5kXIpdGi/FVy6Uz8e5iiuirWd4k20rN0mP/
o1aP0eCOi+2JV2lRglKSPguGym4pjlfWImN9xgY5b1dsNHUYneNmml3LyJvwl3IU
cHcdjjSH10imyIj3wnHp/M+R5+Oyg9TBebJIoIaRGTXs3NDPq5Ph7+jpMkVav1gG
Zqd9UR2rFyjdL6dZevtY3hla9vz1bc+yniJVD2Gy02gOyL8lGRAIwkLYaBr/RphC
pgmGKEKDIPTeuSq9zLN8/ITiQlDxCYeW6cGXLk2Qsyg5bz/o0dV3HWhRLy9+e1CH
CIFrvcbd5ai9sHha9ZqZc6XQFHHJXnqK6KmFh9YL2OOBMr4UX3x/rxr0F7TfNMUU
DzMft6HwxeSNTdtGucr3M3ofUvI2DsfgB9VVr3H3uzi/5nsUtiSvKhw9DDQf3pDm
cF/zQhIXDrgxHHqwGLBEoSY2nlkds1s/5fJU7nkNLzaiiBJpTUENhFBuqz5DIbGt
XprHXNz39E41Qel3NcKJGDQiJVJV4w2aYjiFuV5GQJH6Ydw3on5oHCDT9aQ/uW6T
WAxguXt3ZmdeOjyn5NzkK0/bLSCKbNilXDcSFUSWRFqWtw7Dju5MP2VCGyUZyv6L
wJ63DJ4N4QgYMq16VKB6l2sWw68X0eE6r+1pXb5lxXCQiOHB35l5jelUVhdjh425
Ais9VPLTfedCy8ZM6B+RTUyXVMs/og4Wz5uEbEMYSLHtJVRDG1rCmxOXKVLfRyu+
brBg/dLezQtzUxc397WtjqwtE852+oSudovH0ZqWuaMZ1/w2v6UpaXSIppqn0Q7c
11nX21M2gsWgaLH7vhpoBwM99VZ8E4zFV3X6JU0/GBt0KrzmuHiQ78MuN1KNsqUu
AGlxsHgVXZ7Ww3LuKVMLQdZi995ZdCSUaTAtEY0ERD+TdtZ1mHeJlYT1OIunxjuD
a4YfIXVPpMhtUkptdNvfm5G6p/f5eGTitdqt2ob8lr38bu+fSvK0sCQy2Imj5FZs
xAXvRcyDsRV0Ba/vBHk8X3cCLzLMb0Y6g4OOYJG7g5Z99Wf6l6xXcRfHifMTCLIn
srPR7dBBW9WRrBzy6zly2wsIyet0q+n57lQtXDoJzQCKnY8FV6w33tsIgFZqqZpY
cAt3w02ENJTnCRAx8EUOP9OZMM44oM2FoLs+YnuBh54q/oUQB1OVUx6XJ7q6xbyW
tFv9znvs0rqU+2/PngDZQ/khC6nCE57mrVfnutFfdKxrsrDN1TblzpGrLTeddD9H
e2JT/m3fE4mdL5mJNSrW/CjB0dGmfvGOzZRmMWu3U189UcUbq9iI6awifgrRH2gE
SOfazKbK6ESUw8C9LESS8ZOpgklOUo7nnsEclcFv8qygHutrHgjmdo1XKCtlZhsx
Q6d2Ijl/0Z1su49NIqWExRet+3H06yTm9E0+XI45HD0l2KgChuSxLbvnF4wiYC5T
WE/fCLpFZophYVTvLhtLb60iVSu4Sj97V1D2yU76fAzn2vS+eqmowjFzyeN9ro0k
/6XXBIq73UdoddL/b1H3GwfkunJbABHWzyTXOQakt+xw5Ed3iZQqVS2FH0K+0upF
on7nJ8fQ/wOmzNSEw63gGypxTYONPV0ve/AKfLGLPzKbVoq21knn2jvOmB/TwZlV
EvDRTaKZ70IXylq0y1/tStsBIFiPk/QTqp2/yGMnFP8QXC2FrC20rIPsEGm/IPVW
YBbeXD5mWM4tsTxdcwM4NmZmxeC4UmCL8mlqwOBUP5+Ujb7YiOP7/zUaYoXP5gcs
G1+ZneV0hlMkqsKnbZckmXzgSO2N+dk27RC21c7WAQ98zDTNrsrtaFPdTzemPpP8
m66gIOL6O3oqpx57vgJ0+EqkXAFuwK6IiFYe8ibJ80yMRRNQlGmXPZhtJadzcxt0
cHDY1ng9Em48BktPQCM7oGEVzwFXoOJ3xCNX+oBk7rcJ3fFrRbE4upUfspcqCguk
+umsughWi87+qgsrONuA5wOcYK2oJ2GCrG307p58RX/xiyAEdPzY+WNH+Vills8N
lH++Hr6JGw4ouFOs/xotESkKFQedlD6cQYTGKw+Rs4wHhpoLpd+XOymEKooS6LRL
dmkieJPBe2g7FjKTbhPxRsIHE5ZBGn5Spz4usT4IeIu0HQzo2lm9lgZEXfA6jW76
j3EtKVwZXr6gB8vdVHDN36phvYQCbASY0FGlvyfVGGeBml/Wy9anRUwgKm1B+dLP
iOStVa9w2nJ+juAB6bT1264WpMZc+RnrunHMnGTLNbAJX1sAbYfXtwH2lKdiPX0c
X5qEiuOsXSwqpp3XKvTizT6tzVky6oLiCcUMmuk3xrXxGvbDu+LBYgnfcPU3OwOE
zDX3KudMLe+6ADGOSLT1F/T8FW6WFKnT4tC5hUfbhwOQgfi6MvSL4ip72/VmQT0I
/4N9m2GUmrqqp96KOraUOJ+5vzyKE6yfPMADHr4ohxdQg2itLxEo+noYp9GjqG2f
iRjO2I6BCk8P/nqB14pFUN6ReG+IxbO4i2Ikk2f7KcjJmbDBE9MZS0rrSTVPk27u
9c7KEYKKweXsxNeYLexwZYnGYM5k5mHlN0P5eEoRXo5SMVPl0iTOSnFcYxmX9SdE
Q6P/vB5W1RxLM8fklI3wKIQTEsn+7FJt62KSM7QJoucDeRVS8C7m6JXbiY9MTa3g
F1ESdrXvjoKNhiz4/Re+8C48DV1CIj+Er5Nczcj01p2wG1wEnE5amCflFPvMjn8C
PtfhKg4ZcNF9RuS+7U9O39qhS3p48bUjABgpJWBtWAe94EiuYO+soe8+FP6cC8+S
mqsWt6VDB9/EEmNXI4NJO8uEUgWJgvlNb451UCMhZG2kA3bMn2hAVr6fu8vh2FvU
wzI//lMst2JiCQIMEzh8nSzVG+pjHDFEhO+HaVAjIFtXFY4HWw4wPnre6wP70kXq
8DAPGVzUEdQg/9t/OZ0+auL47hQ7RiEvzz5l2aTHMC0O8FrvavBCOKkAmvhvsvJY
hrg5Ru1hNMKDLx5cjPDmu0sKaPVmFN4JbcGl2c+BVuF14Cg/jEjjp9aSSFc1PmUP
6FPhRi00ya6FOXJOY6WUNX85XlWqsG+GuEbn63J7m44aECaRB/DITJg6a12sZZSL
hpC4dRpMsNHIeRTQsVFqHe/R65GEPz28FYghJwpUBDNJQfHNb/C3iIFnbsvIS7Ij
gqISoWNwUHMvzJUaSX0a+1oritoXUIiPmLlzY//EMkKqsFjBSk3ArAbg0vhtLgTo
BOrBJiOKLqB+B9Z4f353rv7eCn0lV06MpkIbEzAknK9xu/i2PheNLXihdENBCJQS
kO3zZphAEZWSWDlVTua0nDomSWfbyI/1tuvT5Ehes+FO16zRKEOv7LjRztQPHxjW
BR9by+vzdVHFz4ok917EXsb9sBBa3UrU7za+zrE+r5lPBwOtwTbztZa6G6QcnyOe
G96kCywHk0DYAiPfVuDorGdQEH3VWHDNl9xvMIl/ippr8b1ihUx9ojCu9B6AOZe5
OEyFwNjf98Kx91HM8rPh1ljrMemphT4A0IRc8vNKMpjYE1GJnduaR11vP+gRnimy
SUvILc95tz03TeO2+6oVNwuPsxAjUP3/MWw7+ZEelsfhzZZkKWBtioNaFGXP3q8S
R7VxRgHcSh8kfVbkmn4ys7abDEjKJAF2LfKwKLbRxgCfqo7fXuqeRpurePPlyrry
deC8PDyLcyS1JP9OlGZruXMcErnaWpf6WcM53b+I7IvLYUOQfEz034pWkraeiXGl
CpekPgznJC04NZtXycv/eQ6BtECdQnQwMnuoQw83lyDip3fqXk6XOOVl7fzu0hBg
s3jVEjhkkkYoeN4OTnosCXVyqAvGjRtRMVc7m2mmEEYrEeDedkIqEW0PiqJihpsy
cmSKWbu7qpunGiyo+tTTFI/0BY4KVHJl1nr5G47/NhiZtB1BWiMcIJQAIuonGwmb
0a8qvPbCZeTqOv5uHcHCkOA67IujnMQ4eVKiTF46gqrA8rE1Hbr6eW6Kh6Wrf8sX
NEUZ6JkkZRdDswpL+5tnUGa5moh0t1/WdMR9obsEpzpHzi1HNUhU8nnmqq8/8Pu4
XmWuKJZgO5lgKriHQwGgxSSu1u8MBnviKY/caGx0BrmcNsPacb3rF8qTP6bWrTqe
4BqoY2BSHfqZu5/U7OsICgPU9LNclUQNe1Hx45Aag/KPQfIE40IFu+tA2YpzrICH
S+e2AJKofxkiic5xi87QobuMtHcoeVJCAN8qVlb98yIJhYJGquG4JXtuBQvMsH2s
snXdbbaHRdyfI9fCFBeIhurFsvav1Nv8umA7TLV6DPjwiHe/8HyiHg52OIlxpNVh
evgHL/oTxx3Xckizl1J4FJGQqJBi25/SLlS/+rLLhxpo5mcQ7F0ySikGjXCiMrwF
Zw5btUEBzhEpamr0vZmZKzdn77URxRYucNEmeQHN+gZMVIXrnDuCEiHoLy0g0lAS
N/DCkLgkSDJxa0nL9YCG6GlRGgiJYY9eHzcC5JMhzZ0r+g/pVbuHCo11dFaFkJDm
eFqACJWLiU60my5H/ff4CSWCD4P8fNxnV/p+tWUGnRcHUp3HEgz3QiY97G2bKr8j
wfeELpQ04RG+4YxzWGDAcktRtBs2Og+NT5x79WAbFughMQ0KpyqwIS19YmnAdnMp
HrlMJzcUKrYmwNl9Ifn5s0FG4eByEWuOMMppZTtuzNJq6HBF0okNiCQKl+l9Xw31
IdhYLgz+FAOSRaQFzb8nKLxfZgF2tKkysDtoSQMzzo4E/rOWwsI9mG5UUDbUJpfC
Cff0S9gPceu29OVhIBGDeKHo3hg9tpUSA0kPpNvsrdDuNOBfePLyibC5QM7AdEhh
JGGPcE2xVPGGcl0mIC5eCrft2wEsiEf8HaJIv3Il5Qoxx7rScE6Y45nQ3zjTHOdD
MV+rl4StrA6c2n8DWL/xAg1DoBPWSwhbB9Xv4dhyiDK3R1nJoOVIL+6gaqhVC03Q
vYuCHfg7vxlJV5Is+YOjuK+Z3WZD5lNdDwdceimOsJE0kCoaIW7XKS6rmTfvIESS
0NGz7qRj+yRleHFNuLIZJ/1IFlPb+4Qh02t0z8qEPoEVLSRKTEXjTKmDKxaPww8O
hPifZG161vkiIdE/wqrkEsAJNbx4XU6MsoIyYafMj4qFEigfmumEh9MyGeRXqGPj
QHlWTxBgFWAdV2YmndeOL2fH3JPdCwcU9ZSB6v7pXdjZd4MF4mjDbEb0NbJ+A3jg
IQ7ot9iYmfhg32DcRdyZzdLUQaTEHWwOcKURvyMC9mlsHDXHPMYOhkY83T/ayFKU
tQxQ442em6NhIysvLxJZ4WdkaVPfLcrREpk83MILSLYwucJSz2ACsb1UoC9hcuRf
MZipZOVSx9pQIC5x2beF4NzNxoOy0Z1SHN9qvc8z9OBwYtYdee5VLLNh6b/fzGYM
EJm+eX6cIx19tFrNC5LS5k/kFt6TCKXWH58TmDibM0ilm3Bt1udcDSXxHdDoBN89
EQREC9zpyL9dgvWqdq344xFPybBveUnkLUE/Sw9a8J7Pv92BmazU4+SjVeTcHfey
vaALLasuI7PyK4/D4Lk1VY3NrOLLuKYpWMr0he/R0iH1/Eyvi9OkCpFsELgBr90N
d4jj9sLb1IPzIzLUBBs4xTM5q8hnVHcU5bMLwbp9o1bObzXyJLyvaFsrk4KfO5D0
/6B7m/5nffjZv3qHb4xgww0qQi15FX5iKjsIWYsHy1mpkbOJ6z6zzR2olrYkEkW/
rn13hR6DMJ7ngt9mLvtNlxpLD3uRnnkoiT5CAt3fXplJLeEgIRWt0tOOmc+bbqMC
svrbuUwNICqpCyhvciqR1s81Q9vDuJVn8bZ2gnGYYDyWGpDLioUr6RL7db3hCuQW
ulqODZom2O+a+DFpBHlYfkbZo09snEylkMbnA+c9jt4MSxTVak3mZQCTtjJGCy9M
1+DM5EmNQMKQ2BGfoXLCAM9llyuvGsyCexK4dP9oN+aKRlqpReWHiwbNQMOO5i8p
ETUoMSUklqCRdHb1MFCP1Ds6tjpXARyjTfmV/hD0/MVjCt6GflBsRkj5IL1gNW3a
crB7PfN3WYNzhe1dAhsq3iR6K50CEeERHFxwkVEdcZC4OGcPglQvVi60o793eNoJ
EkC3CiRU1U0vGKytQrO9G4BSQsCARkhlDH9DjGg7z4qkp3mcfb9HeKX8EiR7pMAg
0pERE/gRx1188mOUW+LySvgnfKesyXpj9cP8FSAkv5SsXGyPokT8DbKxvWdlI9vu
FrAoZKC3Hnfm1LpMJYO2rccLlvbS0yIPcLikWhDgBpCpEPaB7XVYmSmtbTwh7uuy
TY5VQVeIUthU15mt6xAwYyZqGkWbLuAW6emxD/2se35bTnQWkF+nM1V8nvCEOZs1
blJBkzCeZkuoIIHAe66O2phK4e3/zqBGdv0KlUEt+16WpCdV+jp43/vWaWAj3Ul1
ajNTxqd/GLKsCIrOyzBxKvqsFnnpHm3SHkwootx8CwCJBHMpZHNS3tq3VXo1liBU
qM5HS1UETIozn2h9aQMFHRvrKEXEu7ae+/PuQyPysMSJnGp4J35QYF7/7SSnDLNK
fLkT4WxvOjflbe3m36zN6KLrYUnhFJZ3ml8Rh4CRkO235QVmsZ9VnSf+k6RB7tC8
w8jpzR+TC0HQRJHS6XYf3ZYknE2MLXswjBP74+4G2XvQ9Wc6EXoiM6hjRBAk3IRq
DbURMpNm31bZyqBmAspZDq+dQAnVomG0owT3jODo1xuLNQEv4WD7cl9HKv5hTPBl
H5aNztuJIKsXOL9C+JFu4OTslnqN/GH/7rrfFagtNDVersKYj9Ena0Ffph0lbHkE
LchoX5FoDuAm685wEzMCh/8jPZRgBFNDItjeEEB6MyXoaz/5O7b+rBQ8yoSsa0ES
Q9pRe1fWHwWkuplImZ1jgFHYL2MB0rc8uU+jc+fCtbpyuW6Paxm/VfC2aNze3OsY
6KpCWCv1whPWOhY/BMBHNYnTyi2yeWtZWkLNNUFYijSfs/6G7LwwCoJlvS6Oahj+
DZL0EVMUubTD9VxTVQIhGDDi9J5pYAKeoInIjrA4/bjzvLbvvENKqsk/eee9Psyu
KK0ZnkqfUSGJPMRCd49r+c7Us3A/z847P7kxenkvmldtoQe5I+KQrStatS6MqupU
0JmGQvkaqAwvN4rfPTEVKXKyZa8/pdwf5rxmdjROTtW+0R1jH6ok882vqqWYm0Xl
wY+Qmnc9lerhgwocJSR8tTXuYzBSyR6BZUqHJOc46f7HiMcfB41JAC38xQ1gjjpl
RNXNXRU7P612Z9NHCfAlZ+aMOT1g+V3zuUn1/yGNNEZ8kSjoIDCT/tp/3JzvB+vw
t5725AJXEzwBnmhX8Cktl0BiOdLIDWpZ1UleZnAcSEspdBasmhdLYHTzKak0qKKO
gHLnL4NMqBs/FJJky8FslyBPVHdd/w9ZS0a/DyBrW8IxLnPk4gYkNjPu0bBYzCrY
EGBgyLP0PpLr4Loflx6AzsN81i6CzH7hpQGsZ1H5caYoZzuOgaDk+kI+JP6BS9+x
OTLcjrr8USTiSDpqT/Zcdp9vX59+vpv7q8rLkA35wqDtNqHKQfqSvxvS62vN3JyX
3vQ2tIjlxS2IN2BFkxE2Bt0fEDvO84+X1Oo3o8T+XU87tMvzgdnTXXwLiyYgQsBP
rMr8if0GtU1PgtEwQUA7l5t2HfbZ/L8YTx/ueJBO6FFTXO3i3tzMrgG4eVy4k7H4
J9xfv0vZTbA43vMsE5DjFViTlxfSTWxeoyPeqTayX9rc5TT3HMt+1Jl9oS/2emfC
6aR3WPUlNHUBO2ZY4FD/TudN0h2m7Xw5EMERkXsQTljy3q5/35GxM4/tR6Zi51We
eASrLqFKd7fEIYd/2+tTn8ShJpqi4q32UDdUUirtAoFUsWYipeSYcfSJSoBEPQpJ
IXMNYibZuqCFA3rYGy1SEdE9EitWpdKY/vhCaJk/D1zqot0Dw3EUQPiOZTr8Sk2E
rdZRhTxzcAGfUCFmReEeqQAocedAbQjCZJk6iBupc4AKfsTosyqVupwGxAE80Ssj
4iBs4MgJfYsRLlIEzYXKkuzV51jQPIuEtNTBJP7dGPPZSKetQ6nOdsgoWAEUf3aN
/LvyOGvhm6MlvtbLS37Ej8UAkQDDvxyepOXwN6ZQ6qx2yAAS/ZItjI22zIRk0kGp
HShScW9/mPbBTHe5U0D2ZZUCOvvwW8SyBTX6u+WYWxuUwoBuhid0mNV7YHssg2HJ
QO+O7ZqyLaVgRDrzQFJcPFXRqgzxz8o0tEYzjv2h6SM3Qk4K3VZBevDZchV2sbBe
bSevUKWvBYkUwgYWbcIDSe78Mbnk2I3qLnUCOaUW2k7Ok2gfsOMOWDu1lr7IJXAm
Yn3HVN9dLYNvmqMiBZH/YdBDBejQjxtujf14wsCsxx3oXJggWImSbp/HTlX3T7Qe
bCe8j3FnuECe8jYoNaUMNt1WbgpUoKiovHh1A++5WqQjooxEEF2D/uPIcGpVpjx1
YqVhkaBLMB4vh0RvYXTRaIHz7J5EhV6D16eS46mPqm/1ouXEVee5vxxTpd2nB0I/
R7GXNmdagGLvWbM/Y/IANGnEalZ0Z2trACEu7WPWf61gYh8QXZjap9wxM+vzjmw7
LaKhcJbXJTx3UA7EXlV/fBvBkxv6E6biBwR+5J0G82ShxBTfUHUwuSN+R22sDop/
NnLEwKf/yUZm68cTBLXS8R7GbkiK+9RRtEoWNWgWg9s9BA5Fj1TjjNOUYSMZm4fr
w0FCmUZDjuMEpZYAEIgfoxitnMV8HH/AzXe19yLTA+Ti210M2mgku60itbjvSoYU
8TH2nf6a7/UlAr7/9N+Qj/0O99Mgn7A9giDUPx2o2GuwnxMC757u3ZxXqYrzVitk
IBmqVRF0g0BV1yO2aIBiA7sJP2Cjdg/Id3Ns87okOWOQIYWTrS/lwi6oYvqwILYI
8gCFltDkbWv59NOR/Mmzcgo42OC77YJ7rv5zmOQ4tFBPxwhykkz40kC1nbnZfPMk
aYxoY88QqMDv6t2gdEt6LhhvKWlMDtCS8rF4MI+bt/mVbupXN6Od2qxkc94BdZtN
xE8Zar3KihA8kpCC/rDpx201nyfiC8RAPecQ+km0Nx7pQ4EfFP9AzBd4T6PM6u5f
kaQcYJd59siMzjc/RxNbhoJLPIr1EdgcpmMfQLMDxqPS9hJRThmlyme9QnEYvdyo
rD7j36HaItAoyUqhFXusPMfTgPSWs8/sQZaF6SFnQKpts4qc9tq9kKCUOvQglATJ
Ciq8t52BMhcOeEBxumYqmy53YZV8A6opMqbi5cEnK0oLofPIjp0WjvP+LCpu50CZ
xzKtW6feRKL2l/cGbHU5RjUDgNb9cWAqAKwe8NGHeP4NoNFz6ExQNs1h1KyGM3Bu
+AwPKr+EX3+Dz2qWeXJtJ2uNEwYblv3iCZMQOsMDuz2MKs+0lkrG4X74sNcBVtg1
73EVXX85uzjDZE4APxscjvYsV3GOOEwRjvnyAvhOK43Wi8gpQBoWT8lEBHBmPqJx
DQg5ZSHpRHJfoYYppIZlxdiaXxiTNqsGZ5XHa2h8hRoBrPuofaZdcPJodJbeWUGP
MDLI5IJzKBZMkmqnIEAwpZoPpo3EFXminqgOsw4SDFu5CC5JsFgSPDBoSKw1TZFc
VaZfSLYTQfHky1T4mB5Lqwkr7qEJl68GP6cc692sx/xYXEOShstnSLKNIIwuN6h5
0nPm7/h2d6DImIG3oZ/NsJY8JPkW9GVEe+OLdKNp+D+TRLdI24Q0KHgXhSK/f3Ua
TSqbakRUWF7PylmtIAZvlrzng9hs+6IW9K0vFqe8XtI9yQ7PiGORukmRemJjF1jd
OcoC7pyUbLSM3pk0B52YNnbcgAJJS2gXoU9LAHDHzxIdZF7TKN7wycXTpsTd5YFb
tgEqo0nig9PyyPeDPxJq+Saeo7BkluMxCdCfjhY/7Mzgor05fwf3IEOJHcxZtROt
Rmgrza0ilIyjsvpDbgpHA+rEpGey8+/Dlwgyiisy51ikaRl+5KbAYO0rRZFjDjl6
9FAaO+OHCn1HqWr5yJck4GZ4x4gm/uMYTwMrimJokag0g344OLSbYQCwX3MhD/6e
AhG2LZXweb9lWRiGI/GM6L2KlxQxqK5zJk9hg9Q3RgRl6Y0b5rtqIlrHHQWFwlAP
3KVtWWj5uweRGSyvPAvFGHvDZ2lQ8xSN6RABQzVReKr9B6GFLiiewU5NowD9dQdC
hwTiNWlMyCQeNvmQJF9Qc5QmWL432aOB/jSMjCkc5EQb4Z4iWX3xBTPzbTLYUDw9
8iYpAhwkCfXZrztygsy+c7xg/EpcjT4uUjhQOk9E1GFIPWEJYntCtN709FuisDny
0o7Plffer3wINDXrOWPogHyEjY/oQX9pTt1tPwMh21rxM6/igYWfOsO5t4x7/VWp
u8g4fWKJve0e0c3wIJ3YsQjQqcyaLQLFfhOQ7FW/nsaz0IuaOOYlECChdRxggyiv
d+WLCEIU2mHY8G1SybDH+1BnI3ZysvQI3p+DaF8HRcjlaD4nrx7Wh2Xcgz0GAGQj
mS1WRS9mwXxCWEHKnrFW9UUhumprlN/nrrt1DgS7OullJie0Zf3x7ad0xSnf4J7K
cnyjCnp5R3RoVWPe8wwhqS8mI/ztbTS7lQ7FWe1R1XvVX1CwbjF1j2tKn8gvEX4i
fRDGkTOCQ9p0LsU7scJwJFw2OBpRZkcfVFSk+Vb0tQXfaCL2qfxZPQiMksUjYoVW
DbNz5qVw19fKlRBYQo0RjRWSccBIeG9hq8m6wCJiIbHtUXOpJASwcUV1OG9tUirm
Yo3BCwiByJJUDx+dyNLhleclC5nvPCYe09kWcGeLHPLj9H5fTWnAGVBSlUqAu0MO
tnhY/uc7dkipJISvvwftXC7DzKI+JHVz/0YQUq197YixrJzzequmaPApfSX1nKV8
xKJxzK/cbUvgmoNOqt4DmQEyEvHvObUJsyc4M80qgsyKXB4QPdyahcPYrKR2tsFW
BvvOyGv4V13dZ6SR8kkJEatKPOXCbdB9D94C9xdjJbGJxCsIjdaljqaGTKSWxX9k
tjvnulZcMvSey9C8dIuRzrThQ9hwmhxdAZdACfFaXxBAd85+trNHiBuDxWDCRrMk
KvI3AzLrNlNl31JjkuArAGKa/MQGcrpl53il1vQ2vavDv7HZomY5el+gmsXjNMIU
IZGXFsgSKFtNyQKt+ZhcGrF9fnkH7fgvFkuLpKLYDaNiPCcBt2VQ1aKmXIRBV9Dc
0zclnVI4l/UsFlM8Ky85xQk1jBU+MY5Ysw9xBgbUdqRlGC1tqHDT0GGhoN02ymoa
m0bXjcjcgdux9zkjIANe29EuFohQDiCaRPRONdorOKLer7QOdABRWlVA4lIhBwYu
Po5AILdvcZOYT+AdtTPXks7LA21svnxpS3utFSSpCS2Weh5FKyvCbHeDSIPDRsnN
PpHnbTRwHvi+55CK3tF1MLrXoQgN1RjuMshniJzkUJJkcIy1gs0TGCjpIEOE+Bz/
G/BzK9Ut1ft7Z0LNUkZuQ2zR+ZQspSUiMT8RaDjjt3mp1LIqhXdT56aSYXoQXGHz
k3+tqFValFmr3GGpVjGdcggfbXZ6+jPBk9bqSI2/0rSbeWWaa16Jn1icgq5G4y/9
FLExEuu4Oq71npprtez6Vr6F0RCJsOz1julxN2oeMwKAdDy8laHynTeAmW9IiB2/
HwJAnPfSBp1Z6J61yHRDalMF36kr4xp5z+8ChoNYm4+wmtj8SXnD+KXdJMDnNFtt
WPxJ0fnmq1MJX/uc4/bBldNGxAN4p6DhJXZsx4N7przcRQSwHqdgJ2NYuL44GQZG
h/czu33XKueLZtu/gl7FAalDQHP8pWcXp6YbEaP/W3l1fGzR2DDAwylPkeOquFiE
ykAxSmeqwvWISIJ5cefSmNH+H35Fy+HNVqlXlRoOHr5Hx+3BLp0FLHArkflDWyoD
VnjK4CmWkqq5JxGPL5awyL1125xn8UdbPJj5CJUjPPLFRPIChgxRxA39a4u7DoYS
LeSowHt5Q7w6D7hm9f5KJFyBX7852DNe/tR/eu+3nb52k8mgctKso5s+azrQBp18
g04GDNdCU9fcdttWBpSfBhCQ8ib1DSgHNJWRWWkYD7R/KogRp6aebRwtPgytyJxx
ACV3SlRnPLRV00iMOyFzIdft8CbNvcmlAunyLSZQy3e1GrAbygtT2xz6Jh7QMqZL
O8LE7H81i7HLPOyNAUYjq9K6mTxIAKHXCbhf/mqxczAXBB6tTBb8sqrqU1vmaRHB
vuCSk1qZDVi2T7fGcyfYXjPsRdMes8Oq6Z/ZjpRxK+BHF9VxO/Q/7qesRipjNHLT
jtWHhfty6hKiwpM0fI5dKpndZQA5If2SNf4Y7TgtRMXsl4+2EV8pDbPWQzZ6S57v
lY5M/rYQNluzYZxIa86WcK4AaXsm0uP3X/tzVmRMhE9OumuFCXPfoj5W5rKSd3oj
DCtJHItdZ5iKkBFUAp3Aek2fytHJHg00u3Q6mjIsVOWxjtkXDiyf11oawUlTerp/
RVd2ozRawQPPFJMdeNV4mI7KrbllzTQ6GjOjEOQvtrR/8NLBLlIU7xvcwICGMkYZ
2b+yCaXXugr8VSIXW30/pGDdD6DcSSGhrFKatSkJ73PP7pNbIbH/3mqSuR6vY9VZ
rgjDYiU3xNe9nPZzb4Kdw+QbxOjOmMd6YJbYwna3+AgdBrUfDjJVBofBXK35W8Nv
t1pB3UsSksj0InB+ScbkyRq8A4VsMvJG0VRUyhJDPurRYZ/ZWojLBKt6JcwtZsSE
lUwxon9ykzGIE9MvXXZFWgS8eK7SoUHu+Fgqib79VVahsIV0m/Et5FyVQQ6GlmRz
lBPpb59+77MvJsVjYpMxU5nEyYiR7LE5/v77ni48bF2jDKm7HuG8EAbmtbj8d2uv
JCgxvvcuK5mi8KAmVVP44ft3taDfWrudWBo6qMN1cBYmEnGv35W0IXNMZAgaCxvy
sfJggTz6EAWD39SHOxI3QR/J7lvv8inp8JgHws19MOO1Heh5cFhK/+jowSKzL2K1
NW+G5U72MBPQMDuqptvLGphiN++LVwOWxRPrK/oOzgh7xs7laW7tiABqjhH+dYo8
jnKxXPhM/Jiap91EoJ1FpMjBRibSF+ZB70Ua5bYGeUZYraj6blz1CY8Gf5qUPB/7
l9czxmhuc2/vSW8HcMkGqgDS+8Ae0ysuVuMnYoUvhEO7QRuOfsLY3v7bhDQN6fvy
kPfv/bX/NpOUwH7Hip5n1nmDwLLzc62T8rruTkkLvilk77VtCm6i17Dm0xljxPVH
Khnt+rfGvjt7JmkjCx2fN8oDKhE4y8RQOkrOS9AsnxzKjCZ7k1TMcMyrJp7MtB3Y
aOiZ7v6KKGk/IizqLaDmzf0EQ9MVwHKtsOes3cWnfXNJi+EUoObpSzz2wOBYnoyE
7H1f55Rz3xu39hHn38KUzDc1QwfKCjDz5dD0b5IbPoyqfdW6Dv8wgk9dKifbtaCf
ENW2lzKvXiuooBFhwIkyT9YnaFq1qAcPFMKFQTADxeCpN8MlGQ2J4p/gw5b/zv4v
sOJyXSQaZD5oqSTVTZOmta+4yqOiZPyYQSDD0vLGaCVSsexhTGArv66QenlOpFPN
OANDEe2vO/lbtLQBIVrI6D+MqxkSm/NDUL6r9wsNQoLBlB+a9AaRofgGJTuSfai5
/S/EiwX08LyurMm3Ag1Du88hA0XIcOueVgsY/ujMvQwfIbbXBREf/lyHEGhKDkIc
eCgWz7XoirlHcOiD7bX/YVkoYlRiD6jyomI8xQmTy9mMyWBxu1/8ms4NvOfVhmoH
Ysr8PmM1gHd4ocwdEb8MwkyDUPkuRhvqqmT71L1BLfCP30XsaEjLs2d1cyxRyLKF
hRwCbkpn+DOpnFDnZCS1WcI9IsObs4VWIoomvgOwnckuMt7sd4F7LHDP34wp4OFr
omlZlGADghpvbGFQJJDcnmwD5mpRj8wKKqJGmJjLXM1W1rPXcJh3WdqbQ8tQvfD3
A1y4f65e6LjQmQm3hfLSugzTmjF11BMxL++jWCvWcNMryezlSwMHZUVT2dJA6eGi
MGtpd33U8KnYul/1KH7WM71EolwVTpsk2oizHz/fyl1Fth8mO2ucaZ8JimXzGW6o
8SIdQP5oq/BpH1ghOb1bVwAxjfXUVU5wCZDMz2FAEdcO3XsGRT0jz0bNQrjfcBCe
Uu0/LltsQ0WMZ27lbdFVtT1qkM+FzPV8qGoCx6TBaS86wZVAvYDQef4IRwTYQ8Tg
1c8bQWTkdEKEyAIygcRDYtul3bGnK372UdsjxkRB3LKTocnCDOVc4vbSuN2LQ9wQ
tFIYjsYIm2SFFj/eyHNkzChIcGR2FJKOuL8aFJlOxmUzmTgcX59UfrAR1Ce5MEZ+
IHg3x4CQgbJvLqtSBoqAyKOJtd7IFAeYu3+xuqooBwU6819C1nWevJWHDikUP1TL
zH3eXjSHJp7QKg72tz2K47kw6lAuckNz/lb4cm+IH16DYf40uDEEmCqa+ai0VDO6
X/C3W3nGalptbunM2Cymo5u+m5cxI+pXMhUDNDW1cxQvJnmV7XuO5BYd1Avsiv8d
pfNuFx3yP3/TAx6IdyXAdZALEDbo1i2zBHk7Z2YsXyuabQ9AN/X66ltA3CSce+Dc
WuEy+dwW6DsrdhJGbUxAXE4tKj3SQz5DyGShEZdtBJPjUHFOmULHhJAKFi92qIIk
o6jzzHosYi3gh2WIKYbyjEzjuJU6u1CiAx0P1nJvHvMgnIVK54V2ObyhxPdcwTPL
kAq4xQCOvP3+HQwLSTGkmyEbYrlNEMNOLZ71UFwM4+TJk0updXiCap1iifEAYHdP
RscUmiGoe25T8ygZY9mPHMCTEcVUTh9ZF4XltUfDXzy1d7yJr26/fPrY5DjIUOaM
tOfXMZoeveCpowlK8z79aRv58ZqdK4v/VcwsteKNPJbDXPII4fWUB4ry7mc8PoeQ
1TbpNYT3e+DzEz4+bpfNQEFiKu8wGEIf8vEv/WGUMfcJ/trJiCPknV7Ldo4UXNtq
MQmhgWRa8ODiMjFPBJIkBRhRXcN/jFU9TlK2n+QHBiXuZDyU0zMofR/r8wOxWiQm
vYT0AJMIQqtJ9VXQT+pu6cNqzyzH8tOd5NQezzua5c5UUaysW4pqlFvUHJntYmez
yww8Hb+h657hbTWLpVSMifc5Dpx9Mv9Kw/uxW74o2RXrEljWGqPzTgyFqa+BppFa
nrKQx0u9q5Xm2uxzQoPc5w2IcokK8vf4FInxLHOS2gWOJ8VBvXJ/qobW4/mindbA
mOaaxgj0y0RUu6LwpLDPQ7XjZgHlFVP1ze0hxsza47J6B9NEDz4pESFIQTCoa7TX
YHCf9JaBR6GsEsp4c2lxQHAB29OuPe4pUTpcvl9rzGK5C8RRCxEwo841ArgeOv5L
OA6OYMxpPd1zXbBziCC06GZUjgxbAZCrMJ8mq2jrqH9qS/7wgxdX4thkYn6x8EcW
QKi6FYzS4mbn45NpYDozc7aZQCQv8v1sygNovHW9yFaQV0FZY/oY6GExcrX2auXG
viOa+D0HWYpsy/QCANfR98ZuOcf/PhBDv5jVfbsY4mZvc6P1jRtbS7R1hxyJ3PTJ
zqvECgmADCxsZ+fhV86EhyUxpxokkvQSFw8VM5VevOGsgAMScEm18KpQzvxYmWlQ
mHCrOH1UpNBsZi/T/8Itg8/417fjx/VOWHo1l2BWl8G81IoNnW5r8mdjyyq5jOZO
hEdUtxukVZEnhCsslpPBO2MhJv0Hu2W0ju39sedQq1ETZot1ZFH78yIHLM6qLCR9
oWiL/6q8tXwTf+fjikiWADGqJvmCUlVzB5cAvZyCV5trqg9HDeE972nXS1nDoBsP
yDLcEuQimibuK4lPG9Ew/KZr12+rlXbw2isfSQkbV+Urr880NNkhDJOZ0GUg3714
YhTQP5oY2cycHXvMBeIVI5G889SQzMhCSDumD/R/lDr8ZnBIKGS4bIuUj0IH2tjy
s1/yeL9HoSM2+00WVnY5zG5diYsCeY8unzyN6jgA2oELnseqtFbJxXfOQ+Jpj22O
IeA/GmFNBXBbJSOBWjcJ27Xikw5gP+YEVRSphmQhsULCopAXkYjFLKKFeogNXimF
8RK1qGHaLiS/+HE3Bq1gjaHCeOPd/eC5YsQ1JHkV/9w6jO2BP5k82MXhgcNGjkyD
zcCk+38vn5ZtpF4N8Hg+cnIadM6UFdePd8AUcrBXS8hkgHPUJRI0LHSHzrOmw0oK
yGA5gkqlW2ORVuDvIaZava/tyX4WbCI5j9lylfLBArfQAjnOOaRCxoS5eMXHluoV
BkcCPSLENvyMl+9BzUHrj0wytROi0nFeUd/x/rdXYoamLK67pQgPMJsgDS2/eKy+
GwXNTfgIOz9CNDI1wHW7mN+ehK6p4vXCWEoqrOAYtEKjI/IML8rEqYlG1vToiUdR
n+xYcs/0Mqalo8nXceBbCAqioQUYi/Apyl+qGIkjRJhhWvBp+GcSNkZa1zsrh7fD
+qNxibSv/OpsNebbyTF7p4pmZKbrJOJ05tFG+eTvmUnsPMt45130RYTP2Clo1om6
tD8jRjT9cV35wlEOtMYW0ohbbGvrZbRGQAb8E7Wr1cMssDUA/xOwfd4jUeBNH05i
riXptvU0xzAqlGavjTUH6hdcTndOMH99bFsiueXl05uN15b4HaCrdYe2MWAnw4RZ
fFVHJFCGJOa+KBYFWdZOjPsgCOQauCemxIyHRGNRyGQJCSeRzBbeUsxZojf+cj9r
xyV9XbL7zOe/MqrnQJv5TKUVrk+ac2l6sVB+oGprmvFvTeejy6Rz1ynEMfbzj5Kg
991h+RTtja7k+5m9+hWDWD2GD7SFnIuKUMtcdAzbI/vfEOue+wTknCRy/zKixO1L
AovwzVFR34Du8zDmfB6lnzeWuxirn2ftZicKOB4mdL/XgQWkrXGP5TO3ZCgw19sp
Ry/WNy4BcrjXfuIhk4wgNpHwkMeQ/avNr8H1h6nBI9NdsrmyH/0ch0ACgQAKGhFQ
rrvQZO4+aNpgTKgdAIaswCc95D3rIyI1VGKdCFB7pMDiR9Nb2vB6kKuuyv9iJdav
E72NCBYRLi6PIGGwWKI2lSqoGtoglFhLbMDsJoD3yjazSHWfhZGRaapDvLZ3mx0f
VU+u6V2WHCjOY9dOdaErveZsdCHGn2+QefJcBY89m3X7R9dQnp9CQJkbNR+vtlLQ
EwBenDo6/gmNQ0zjjXWIjaVfya3ugVEZDzXr7hx+R+VrxGRimf1HEfaw9dJRfw+5
7wkI2NVeRdGOoDXiTOFHrSyEThz11KLij/HDJSb6i2KiDMt1fQE4tdWFCrJhK3Lv
P4A0SK5bVW52JDaCEetdOkPHuR84CvE0twWgVGOleEbK2PXd+9PZS9lMg4k10leJ
uMXIL7SMixYfga1miR7oNI5AusnTggfQZ+h/OJRK40KJm+Emp8zIz1eD96UQ0Cm+
0fduDpeBXTLtHaY3DFRFg1GtEy0w561/cEuPFf0ZoczSHGKdGyBJxm3ehcIh8eB2
/DqLca45WOPFrsjq+CNsbeT7Gp8NGSO++/hPKGFYlLAbQcEf2gfSj2TkGEstcwkO
qG8VgJc1ht+WPHjDNTJPUH2fB7ntgaD4VA/uuL+S9pInxgk+6u1s79rvsinLrIee
/w8rFWwPbre1drw50nIFRaR6NmUjVDBn8l1t7voNGmQz5h2w5B7okMjKUmfDdi/7
/X066JcfIL6wNYkFm8VHFAH7bCxC1oBm/gnrdrUvsVJV7nQxW3d7cIWL6ar5iOL/
txnU3MWzvPHab7s1NnAPXbiu+Sz73wFMxGCuc9sza4qOMsE+VYc/fi9Hsfmz+UFc
u95I+evOhzSX7hKfCqCiU/Ojum+i9610Gd+cjORYvjhYWOwt/MVpadiewOb/TN0B
ZTYeQzqGEl8soLUG9hipdWXoUvBSiW9k8DHQ14Illl8Ku1kQbobVCyw3xoUtaitL
iLhpzcf6Wv2aNNRi15NbraWXtaJyhyYn/ZCwGHP3QZE0hUEU/GWAn3p7+6jF7Whl
Oq+8v38KiFZdekKnDqr4Dt5+PndE7hrs1rfoTzM/w56qbZDHk1tN5A2WX2r70qmH
P6yYkb4DiATjMLplY0bFKaaClv5WWVg5CQCcTfFxeXZSZjjFzoHixZ96UfBDJHlq
hoq84YTAYN+cYwvLdkZsIf23mXz7pSLPWfDjcICWZJdTKbCqI8scma9Ra/WqSuS8
hiN+w4tA+4GV2DIcW4XQdi/nCzXaKbcKGBIy7SINYJ6CthHCAa3L2xz0Mi6J6/Ae
Ge/ivofSCTxeVE9j61ZC8P9D2F8M+HCEyLSZHoRmridPYjkiHI6sYe5IOBAn38pL
XFG7j37bQy5oxXNberVqGq+DEnUs5C0CWhyVyGcgzf4dqlBa0HZ2l/ENPaupo+DG
hVmSaqrYES1Yjr/WrnR0f0/wCnM9cDfeoY2Bu6KF5x/p9W/3KsaqwSfEqX2D/AKN
JGugA3vRQTGBcwb/F7ZHpRXKJVcEHtwvAz7VcETFuwg4kHZ/RGgR3jXbPOtm2tZ1
RSERCVteE3tyhu1xhZ8HsqxWtuEjyrjdGIG1fvBljtPfTWmb4xf8fawXPcsDSbHx
vdp44nxA8PNwQzKdUVKv+7BS5V6t8neTMI2YmQZhoYCFIAdGw8YH2BRreVJ/P91J
4GRw/vIzRtKzT/8i9fDtjbdut9+7G1uIx53DopVSumsqvdEHewbCkIgPvHgJQyTP
5FDdJM6AJCiA0Zb812lpSEfJavvMNT+4OnRQiOtNehW/PSyS0zB6ae0YyUp3kOBb
Ta0CEEXIymD8Aq4Gzka6sJ/ESKF4J6bVVAFMLYKqq5vA+feBezGYwFsJ8prkmwqZ
RYyOVdA7zPRI6qDg+JUgMbo/bVL2fiZdH8zQw4RxYLg73XgLB8mxQHDr3bCs3ZCx
CzL79MLusyDAS/qDOYwkCAPiJ6m4FG2kGP8KDejCl39/r5tC6IPsnEQJjR5yKmdp
dwCmwVcKbqRwUVvXEzTmVNFJiG4MAHr7/D1ERQEwWgHMXXh6XJadOLXSWMM5JofV
+rJy9Po6b7qWEp5NA+pjEPa9ldTJ1Dpxa/vIQ0V7Vgdc98vT6/8B+nMQ4rYu5UeB
NgnvWgBYspb0gF8RYE3Aw0Lk0z6hYWNbRO+xj2u7e+K9fF8eyYMjiehjo8TX0Ad1
DEBwD2XJFs6ceQ6JBg0zG83KR42Q0L+2xDrALOuePZFeTSJEgbGYi7MXZXkQyrsc
uF20wdSvZErpIPnP8JowNrh8PhJWDeeq0XtlYjw+cVENNvTD76xr5GvHBAT9sgVq
csSDOiFOPjB5UFMAzcHo5AAN/WEhBN+5Fqvm4Md5bBYsBCe6Evk0VvE7axOEfzVt
ansfh9hKvWIi/7dglj0uYapg4tXZuk705DSQCsMLeBREYDsSW4hMGYxmmUFvPwY+
OVt+dazpl3CTWYpow2tFqHOCmO6AUlzuy2hwCTYlLSTMpHlCB5t2jfo9zIoOfq6h
HOWuqlsrNI8PSCb2xhZL6n+j+M9GL+gabStIcKZmV7X7x9cCxbhGbvrCzrbakd/V
L3unw6Ics2uDIgRyJ9gG39zDNFvbwX/zmx3WOUPug9UYap+EJHQXf6fxjEHsn0AB
FCyx2xUox1nwRr2LmAHrzX6WvPh0gn2bNn+AuKYjjYWA2UA8Kk0yxSBfB5orKNNT
sZl6nGsbR6qzZBsotj8eKeK052xgKlY9YqQJ4LSgG2tadZH6zpReUAiHTg9eW1yl
XznBME2ZMC1gZhnvM26Xw1LxXFfakahV9rkI0mRzleAJWJ55leW1OwfoEFb9k8KW
Qv/c8e4T/qIreZkFoowBOp76KcQug5LEiU06uxzgnX1o07JStI8XUfGteGtnXZDX
xo25cOrEAD+iZqM7DERI0TgiTlw7XgahBQWQZBd1rJ8yhGB9QFbYqvs8LN8HjmKk
hXJbch1DcqKLlXBAdGLKsHOis6GGPQsOEIz32Uy30zUfmlt14geR9u797GVUtSuW
mkdge+ZHldy4loFhT41uotOyIc5NKJpDUp+BF0qvIC5NV0Z6j9rSV+cRMYqcs9X3
UZK1kWhrQfwlD9npbuV478OHmk2ubYuWDGAmqhCf7+s52oaEfCkUhT3OtNkAHJPi
14Ei9LdfSq/dTxRD6Li5HI1d8J+K+2YkQzG2k1M2GlHB+c84GSHJ2dmBR7YfCXDg
fZiXMbv9AlY9E+m6EVEwuTNoW2Sc9aUUQUuPHeNcB/hQEu4J78AIiQkqNX2AllSK
LU8Mze5JAeIdG2CpmjoA5FeDDQNg877vK+EkzSaV2KWjsxh5AmYnkDssqO7Y9e5Y
Zs1D8L2YlG5M1u0xtPurfFouQJlnCuSRQlUhZ0Is58PQA4kkKHNr7R49s2z3PBl+
FDvIARKUXAsD7UaJGUoemOwX+ouJfxAR1IFxzocR6ZoLPh6MIrDoh6/bDw08gdYY
OoIcKedlFeEoWaznV7cYEBiKonfl8sEr7y/tpsxu+GgEQUo8ZM0kSdLIxZfyNwjU
gPM2AaBY+bYOvK4ghd1u70XWuxPS26rnSDlsmJZjzo9iR+GSmZSceJGToynuOs/D
/w6dxVcDy5X29SfLzkSzf6cKsoyuCpx9jeN9LppQTIBB11O/npN3NZqKmLz6nA8T
Hf6BpoSpoaH9FAT/H6KjGJs4VIi1HyVXKsip3v+qCQhM3fFiva93KGCTjXTWurTi
K4wXW71lKQLGKZu7oBZaRBUc/1z/UN8Cm7Z+Y6VYITehfXp6gQTIvq8gBch5Pb3n
c8DO0LstaDqbpQr1HHWvJvZYW1vdJ51xrrVMcdsS8pMg39vq5eqwaU5Js4ICO/Sf
5UR+PzUDTV6nDWBbaQWSMC95NKjWJzjc0aJEFHunOPaaue28wUBpiWlxFGM94/oC
bt5V9rEKTSBjFPFq6w36kIx+ocB1DwPIQVR4ob5WnclycLcYaEz6O+Tij3JNK4iK
oRK4Xi1hLEHJjL7ab7X1mQSPmRKm9arbyRXrnCpWwgNBe1h5QT6JZRxDH6kpEmmO
DCtbINoNmMHq15X8B3sr5Ct5Qr33NIaM12eGbjsEJzEx++G2u1g/unCcuJNnRk53
oHuEmusqmCiY1ouXPgvcIKum40cGQYWKpUkQ1ePBIkWe8QT7ryV/cndHHbsUqkUn
brMDJHyJ4f7U3GIZN5o5petO6WaVMEdjaZ7TYMs1lwy2zykpsWag/wjtAe6dsA+v
RjnmwShcIhmNt3slNaguRMwFtcHXVqljWRB8ZOJ8W9DJm+Cssb/SFhIpBoxZEN7g
P31iAbATcXl6Quhzj1JFcRLiV6ijyG0Rcg2f0ZVQgQ0z+rHaFN2mAeOrfcA6Wieu
NLZfeCTZtOsqPxa250TQxdhVKOOrEPywA8CpDVT+tH8RLkxxjtPwMpxo4UOx97fO
sYx3xCFEnvDAtoWphOT2kWEZJXAlLfwX5nW6WN0bt/E3Uexm06zbVlpCANq6hpCx
5FjjLMcxumoDAwoaS7ukjIH14pCW8qHln2NuyA9/yGDuYy1tlyfIQiJWR15kHVoY
p8ZtoU+Iwl1B3my0vpOfxgAfhn0Rx9qvbjRmaClcMfJngwvl3NrRufCWy06WEEN/
rWij/SnDytiDfeQmhI0NmoluRBEQMJosTDvxA19RbyWMeM5ULAARfVVq19d2H6/k
iZHVntFisdynq5h2VkhGIlf3wJNFR1cLuLj8rPQwq4xSPi/xrwCZNRTMdS0IpKsx
fnpTJlYVeEi5obbqWheuKqhrVuRFuC1N0VkTHL5ywkEhjPS00091UBwT5Ch7OriO
Y5nMiTw75X+DW7QCeYE2nQrAaDe8u9qYny7bxmHAG2UypN0HluShkuhLnNvwd/Zg
fbDHI4JEnr/PBhwP78Rg3D3KBCUx+KoANf1aZIOYYq5gRkl95BeHjIpzekYKPaY5
KT8IlxaRltBQLoHP09xkFajae5+56mzQSv5rmmcWA0Yj/LTLs6plVOa+SYh0Yw6u
WtkqAjz+HnKF6Tk1WEMT5kgqEBX3xAIwfmY0zXwPoQ+f1KP9cj0MWBszRU2I4RrD
baVdZE8AZva6/mc0i/XptwD5kBYSp1eLHxCS9NvhDUFQgVCpekh9o/SfWNPl4nIp
irAdHf28wLZmi9NRzDuZRBKAhT94op5NSvGh8hQ4hHexObVVoF69xYjJ1rsAEAL4
igxLUSwkHPZ/6yqBOGzgGIUVTxuihgqTvx6n6cF9Co0Ik+Qm3plSuS9XQLY2yEh+
4eEUQaJ2/iUfY726XCxOVcrHjmmHN0bi/p646F9UoUkVX5vq67O26xa14fRgRZ8e
LI9zMPXHPHlHDE95iT9XPAZgapBBH9wbmk4xlPdop24U1cK30ekxteeJtUe3y6Co
wk8Q+2yfJMypiJW7JWafUKnfQktbZXaY0ZYwbXbiaZWMekBFQ7uO8AH58O4kgWiL
mZloFz4UoX863YzUW/alVXFHsxooTLBX1FKkuotqMq8OlDh33y4/9OxNyQsmOLXG
HUY1p4f0VZVpNdrPyC42EOtEC6atILYM3Zk1K97sO0kTV3GYS1IKUT7cwN2l9Xh3
CsdZZEJLwDMAqRoH0eQdkXAgxppHJPMfufVBy9KFWao8Q88naEMVmxiwMPfFIDKO
ZB7eCIvUd0n4QtVjnLVPqCODSemG7NWsqNIzm3XKpkshYyG7nrSwf1G2QY5eXwSO
HiWvvnWBPXYHsck5jZ46K2WZZqeLRBmfD8PvWf/f7ktQCsaiatr5A1ExoDATrXfh
qE+XxIqCmnOdvD9HMw/Bj56/rAxPE1ZT/NXVb57ynHnN35NpoTDA4MdgsFNB5V6b
No0N4UfnJqKHEk5rNOdPB9qkraVY5hhGuhv2AJ34JVh5VLi9nAfLVTmUZI3Hxb8T
/0IQQBCN1Hh9htHrudoQb0RpX3uPt/Zu66g5lHbwpx7y+CnqckXCWeAs3ULX822q
bAOSKhXivHWgRfLTTux+QJPJbBjhoy+/71/7Xlwu8VgfGlEXzabTS/wbjMjyjX0G
DG/LFKK8A9NHFF+Bh8+Ez47dGDtz5XLVg9eYhfymSbfOp5701aTKDoYqt97j2t8+
dfzIsQ4xIXI+xq81IqTQB8mBnOwXbx3zT1N7q+5F5lNZZW8t38WY7Arp7ZT0zzhX
75xPZtfNQnDyxE6x0gWO3ele/bPwcf+KsKsDOHYUeOvDWFhffI8DowIcqFSuwTp4
Awt/9b6Po1TyGRfO1Vvogx0RdTmNXucllsD9olhBRn4sTvI8Fk84O/i53BPdr6ey
xUox3tkfyT6CQt5uMJBbHuR7SuSlE0E6tZRC2+8Nv817j+xLzk9L208hPnedARRZ
RkB5+acw3XIPsJSmNbVOjrcFOpLd+ZXRl7OE1xN1bSAngez+VlEQHoxld0a0omvn
dsHr8txeWwP3WKVoSWv0fh6vM7u3jKYtnnjWsf2/rQUJ+eZ+HMnFq6XODLCLo+5x
07paa8/DF0V/CRBqBogyrx3wadF1tsmJABit2upJNrQ1buttKH3iFfXjEwCdLJby
GWUS73ph0XY6YuaJal3pMJKgrjkXmNh6+696wGUuj5+bsAv/PsL/un81XZlXNruk
YBOU9q5pCT+wmdwhqKpcr3PxOKmGlhW/FFUFh/J4BGh+93aiNLIODaZidQlDqA/H
u02Ni3EHgwM3njIYEhCx8zONFjypTbNy5eS2BkpNZgqLzaBjBdflwaMk+Rv/D6Vu
3wA5NAIYVVOYlZ60denCrNuYeMaf9RMzRNtMluPz8u7fvWVM0sAqr6Ew7/FAkMaE
8nMZrT/aFWmPWYIQyNcpu7hD6/kbiP9qjcIBKcl0kOqzvQAAEGHbb2oy7CKomaIB
QC5BIJjKdRhwH3RF8yaJ65cgCi3X33Z/LwfxR1tjBDFhPrW6GEblIWjukx0koO42
y44Oha4WUYK40Bah9+BTjTTdNK/V2hfAeR9LPybdaTKxrXZBLCtvmujfHThzNI+5
UiCUrPkl1jAGnGnkN3kla0l9PNhsSfU26mLhEaEGdBTYn0G9P4zCYXzZxTSJuqef
OvHyTYoLPXbuo+hOd/GiSeDI2UIqWZ/LwrvbY09ZzW6Y2y/vYt+BZHim4evWwQ+s
HFyII4O68zyTPPiqCuwE8n2MrB0h96/PIGcZn9LvF6CAYLT761NbO7JjAYnIqKOf
wfIOUS5+JDK/PeoAG1sG1vBmkVy9m3/5eTAWCFZbHABENLUZblHfUzJJDQuFQolw
zblCt825/a7JgEP4HVcN3GCwpmIsGnnkUhXVkXjFvFFO6s2BgjEBcsi2iSnMZ3VN
WaH/MU5iMeG6d56X0WDOJOUXtYfk0ENFDn9GIuYC0MOPhysCVHIgFYe11nMfVAdQ
D0akIJkaLT+mKEEzzXeNH7SPcajrzWvq9mrtFaGQuZx/rPONPRMsKbT9slKhP4/+
umFy/psutp53q0oKedm0pRDi5KaaWdwCKVYTETkWAbZUuSEopY50NlmB1GyOfySU
AXDV9Lzs7Ijm4oN/CV6stznR0Z1YtvO/LkXBYiQwTHh1QgGuCdtlDPvONV1vW1JU
zgb/5piwy2DZM40xFANgp9X+0CiYQQm7TZroPsfmUk7fjHJZyBxHRFOXY1Q27DeG
l/Vcixd28QCqyzmjdcrDtZQ//pkovyxUNwFNpP5kx+T7d1z5nGgZt+XLYjYriDz5
UFlhUhU8GwssIS/TjWteggDwaQmdowWxXW0aYZ+Yppx0eusCuZb91DQ3yz/FP2V9
/tk1KfHT9dAHfGy0Xd8M+daJPhW9IuK9AXeOsGXZ0h3N5OlXwmLYONXCBVmxXoA2
RGshnlRJ2RLf8q/AMxbb37JR7357aKyHZhbbm4T1YjxrGAMXRN1E/COB07WNxqiF
QzOuj3FqySmwQZhG3ROBE25g8Jt3vXtlFUjF9FIcTb5q3D+jJCH+oUP+dH4dqD/G
bwa2Xxq0zJdVY46inejJCSlkiazU6sq1iWmsaL6MW9Cwct+sI//Uy90KNG72Q2gL
Nywj8zJSDRe5v/90T8BQHrhe6pLREZSdsB8CJwstptvmMnbD1ZIZU5ArI1CS/41c
mmvTbsW1etr8ZQo25ea9HdS/E+/GgZ3KNfqoPHH0bvRBSYJ4SNO7WQuwtI0iAZMT
NE8GkeO/kcH376bQ/dNOy5IPBDrCtAN43BwB70OuyMnQjJDDdhF9OkV5tFIhdiG/
eQ7Q2lX7RplGcmEK3wNXYJ1Kj+QF0NdxkAopI97OdaIZWeC3o/UQSI4faTIgPDHI
/9Se0UDCe9y30PxESs8e8S2kSCPhN0DEL6Uun8sFCwCV4Xn3zzaJn+QLtaLdyWcF
1pyRO2xbep4ne3LHQvf2EG0377zvXCyFkpBj+GmWHODLEJpZRAvoKfduXq36frUW
5gzlMJvDy54QwwiRvcfw3RL80iWP/45is/QEoTmr8TAiQR+4ykv8DcIqThRWsMtG
XslHPbifYBbCf7HdIqTY4NXoKfwCaWcqhOK86yLdSxuPuF90rZBgTzjum7Sbjt51
GhtHwR+tuZTyurboodOFuT7k8xc4WMZfPMU6FKt19xfYYs0zSU3W6Ohe/eztFKEC
EzQsqYJDu+uGJloLuZPcWpy4uX4ahNwj3vKg/zqD8Z0vw8+mTwR1jkEwV0gxZc7n
BUcFxG877Vvgv/4bIPXiTMWi845Ui7qfsvmxGFj7YzwyhRnz5PoQ8hib+Jiy5m9Q
eqQh9PalUlCzf0hMqhGGxNgFAWqA29rIfPrn5ictIS40Q03ToTpPzEjGsoxRT5A5
K7bHUNM7aaZx1eCufG8my6FOHpZAiiiF769SlUD50cNocnE/1VFNPpwlBYYp7fxn
TSGVSjSzcGIV+88148ikI0oaAezfXWhP3S8wy/BVTJjIdE9SvvRseHZ5cIYCpSI2
p4Q+BGD+wK48NBc/9uMjgVuRJd+zhlJe/wUQoofAJEZFq48hfkyO0RdHQUWlEP+w
cvM6vUNbxjV4u3L2pxCWlCYmSXqJHEu2x89hOrIXShnxfz2NFEGJsPTd3xPIKaM1
fqYp9JcrSl/1KQEU/1MnI5uBs3e2PwCV++wn+fdYQXMHQXvPnXIyhfu3k6zXEj4C
Ade5bd3OdtzjZT+wHYa2z9L7NDMWHN1bJJdwEOcKTJy4rRC97EsaGZPySprryGqD
LSFI7OUCY520++xJzCMTFspwQNtVBWlPUC1rdAnRfhrETzbldPjsIo5Fo//RKRtv
CRy3JwerPfP+TqQ6uo/xoe02Hes/vNr/wF74o72yetDIJ6hNnmW8KzTQGgK++Q2D
wPbZ3gJyadrPdkqeaLszVAi/xCsRY2rqjiapyTB0Au90fXi41U9YYNIoTW3Kh7y1
powzUwGAcsV0W8Qv9+yoU1y7H4xFMEJZ9J9ao2VT5c61lGNCprXjEwfvQyk1Wjmc
ODmvLKSjj8jMzH6MbX+6iAsKuVWbodLNsBq4ZQWSDcNYkTHTH8oFdM1CqB6G5ey4
UnATIrymcmMZbYFmuRekXgpNpieXfPXUdAHYgdeW+OsrVkcTykgaR4+k9eEAXKgr
TiU+W7K+ETWkVEqOdMlRbvnNwMeBafhofS7clfgInG8Kp3kjUnnz7g/RCa9Yj9XB
e+Kj/T8F8EAmk8W+vnltjS3u3xvGYoi5yFa/LKVlxU+21/aLCoE7y+51bFnJfqQO
Mi0nX5IGuEqUUyiFVC9q4Db7p0Uj3YUD39Nb740r6JtLRuEe3B2Ny4mwFQFuzwJJ
tPWq5IBLFPs+Fz9fNViX5mE2HaSV5DJvAWNZ46UbcqtYEoKyYEwVmuyQdZ+3CHa2
QkZlJ2gXbf2u7jW1UB22R6Di1/ub3mM78UgXhA6Xr172YcUjUwblJah9TvXcVCIo
BoLcJ88l/OeB9YBxRK0f4CqviRPhMcLfq2a/+u6v7fj6h7nqGWbpZOpGe7J1rg/n
s6srWp7Asu7FGKAWuzeul9yZL2sXapHUZSwLwZiHacc97ZYs6EjZUR7/C9dqfmDi
t59LUE5hwsds0zHDDxWHZHFe0P1T7ToX7mu9ObPbOAflLuQwd8aHXq39ea2xSGSe
XHdNeexb7lJ2str1Gg/bEfJ1fm+3dTDGtnkK46HS9S9LGRE6AD9jZK+dC1QH/xjY
AHV7Lv3/ZiL7voOyChF8nstdFgnlITx5UbUyhJNCx++FUnZpAQP03mKFYBFz8yZv
khk4b54caRH6IOADIq5IIWPCvRWAnX3ubESp5RrWfWux/2zml2sRvib+Mh+FIuCh
UX/D7JOik7k/tvFv3vmMO7MftmhFM64/KEaCQtHyOzZIN2KBXLJUp7VFo7mhbViI
Cq+yvinT6dNCBEJTNW0eNellaFANEw45jJjlAu34Mk6G4AByJokQxQfWvh0TLFE8
EAMffK2b/CHHEFgJf39KEOcqr64N6GK3v+ANmc0Lkq+USw5Koa9Lv4uUvpX89zdS
K+RQb94llQFfVEUY9qSuG4k9hg+HNVbPOruLvtr+1Ml4UUvp2uWprZdni0HiiW5a
KbhijY4/qzLEFuUN8aZkj50JwTQhP7eNjjDJOXSm1Fd0kEJ+onU/+igP3M2KlCzG
zjInjef0GvtZ2l9BKZuFhtg6tQLSNtVsyXO5ZZJ506vN8sMvPh/N0uPF+p5/wUQM
NWzOMLgodLyBVNW5wystOxH76R0O8K6D2gbAVaY5akCjNINfFxfVk3zBw6Y+mldK
cZkpQmDA9JXCILu3sCHlu5EgfOGk4iRyISG2+KVA19c8QfSAy4RvDEc0LBKYfWZF
7E7AknW9bO5CnezfjJP84U5sOVDESGpgvjDs9y4tDY1Dk/jXxgSq4zuNIVifxBWd
474NZ/4/CDmdbZixGYrhRJN75QTjEm2Zr308dTwMPm9nN3khR7TnTxmpyi7KBBtA
/CExSpYPPBRUtPCH14RCl5o1Fu4tF0WCZ8AARTCxfm6SICuXJLFKLiCCxHW/fxQY
CkrPl38BHgvZ6EHfDkou40YddefkWpclWR6PWducePtjxe/6umYIodKw+aXW1YLU
IcQlUGQ7XJXW+AWGmJ14MjUsQrCpXKZxPH1ARsGrCBw+4xpUYlkjMgAxwGi6bg++
S7bZ+MaFaOx1fD07mmOG4u7YWpmbIFxvzJJuQhnteHz6DKYuhjPokIpyKL3PEgxb
yshgYhd/0f5Z5GqXraS+F0nTiG1twjrBibn3HCW/UoVhEM88Pb1G3ZzWGUhIkKvm
x2azT6tKfc0wiFdv/QfQ0BZvZg6C2daEPl8aE86O/BfahkkSLE/uu8CTT00wtWwb
H9LJJIuwS6qaDapyI9rRCZqkfFmM2YH2ctrOMm74jbVR4SC4P00HNaVVX3B8E6JJ
Z4lbhtswVoRObDRBSYwzTG8wd6W8AUMBMHc+hBAg5W4Vk114wXzw2J8xwQjIfAd2
mpWXbdbYy53Dp2+HVvq5drxNU5nbUZQXB2tnkkozLT+KcMaNYfqC7ybKFfxs+igj
P+m56GM2dRbDZHdDMfHn0WNwv4fok8P5qsuWnIzN6SMxNFlWA5LoIXHObKNNsPkm
mbwCf76+1dJeontr9NAG2m4FKbft3DZfy+SNCXF++XWeXB4yxB44hZRMnF57kreQ
sSe548UGw4Sqm6JvIjnDxdJiJFMAgGwQIHoaS09SOnfXglqQ0y8yofJ8qube9JjN
4znV/bM1jRpSXSsFX+sh5DE+zh4Wq7bOf60skgWroHT0P8XxBZm2jtRmLVvY0XoZ
AVV51MrfHRkuEhYmcj3O3fvC0cX8AC8QTlAUms8Qk8nJ1ETBfSElPlFdIwuaaO39
KoU0YN0DUbS844pPpPwKD29k9j8RAHQOeokUd6jT3dzy7P1Ht142t+ws2bLycEa/
Vndcklgy5UXFOuw/DUBhX1XJBQa1IKlbY7FfxkmX4gF15Y1pnYM5Ehh6KccWEkDb
uDiEfAX5eRxnMOGLK7sX6eSNVj0rhs8aBa/4mGW+tludEdCJIiZ/jnzEY7tBOEu0
X5joIBubsJmWI1bCPtPMLRODFcQ3P8ZKnS4dEP0nHYURZJW6Y3hQiVtnDVVx+ojV
bDPjHyJlQqeTltV10zD7nExRTNA1LVnp0154Jt8dgYTrxfiXjq4I9vquqS0N5Kju
dHdvln6V/V5I0ByHmVfX8CWxrLMKtKBSwYNhZARw8/gWdjQl8P9yr57vzMlaK4kF
5+G7+724/79OD866uiDWzjiMSk6fQdMbLeKtq6QAJJOuBSGNIXdJzYFvCcckjDc8
jJUiP/w1538Ae58CAnyFqse1h0gr1P+OUdm0B5t2jOGRo6Xy8B/TOyiYK92FGHac
zFIl0BfP1a6NKYuOAtzb51KpkuydV2FIio2qEsTGQCoH740n33Q3vUGysHllonYS
Oufc6ox5YJcSiWrnVMRXE5Uxq3yTosOIm5WkXLU73NsLphGRpe3HiywVV1ll9KqB
8drKI04ew9xhZsQfkYOG+uqMryNtS+zX/3kp/RofISPZ8S48R47z8TuCjBmzJa/f
GbCahN2yU29laHb8YxU3fR+UAxaKifzL9j3vxKxhech+VM6VNTU3lJfCnXO/z6CU
A/RPhCe3wF8F8MaPLI4aYX4NNhBdWOlywCaR1g32MJdXFIsAPjvTFgjmDT+NpU6f
EiYXSHeL3FLof8bSFa54QLl3/tvdu0hVhbIuZm0xikDd8KVtRQyLNUxptpzQ1+Yb
wV5EvUJlungVa98UrRKUrg6STUKDMH9+2ag8k7RtDfaeAR+698Nv4zPKZ9TC0QYS
Ejo6XnXzLlZa867NNsh23eCUzuUeFJdn+5SEAyqKldRclTKpFgqyLuvucOm3rr6I
jj2ZrdCZz6l+Cd4Zllk+jH5sSvKFyV3YVlE52e2A3PVf9gzrfvQZutlgYaAjUt+2
P3NY858N0S5bykxlgJ8JAMvQcO/yRvGkGvKllB6pzKTsPYeSlxNNMICTaDXNyKNE
RxPq7U87fqLWoekicKaEx7uX3xggHzaUIiY7vj8FKP7GRVSci9WzNQpZD1DngnOk
1aMNvOXRp4ILxi6+VHT8qtCWH4NJY60fdEkXllta+SbQ/UNyAO7BAyD1K6AB0vQh
z7pnstpu6xV2xIfnv6oeuALWTc+TOVsc9fK3nny31Ul5xdpkdztyQ4BQtlTnBbgY
PLganNPMVcaUWaXVTRtC0svcJ//tEoJh6L+Y36TX2+0ZOHQiRwtt2sVd4RM1ObzQ
/tKc30HXKXMXBNkxLls4wqXD4bvceG2+HZp/KFTfN9sHsftTL/QRjGVx5Wa1BTfO
MDn+E0Gl/osUeEceQ8QmltSaR7AGlpyWTV1rTjTD3qM6aqFXzmAn7bRU9NhWAdsq
cxjXxTC671p9soVXrCA1wEokhonM7SW5ccoMe451bulVzMiYrECTa2O+IKpVBQ9V
dlGlBao7WNBD6qwgoR80eooIYgBtSig3ZRF1lHNfJTqPgLtP6L29Ea2YakOqBgb6
FIN5CZT1Ga2CQcFF8G87T3OYYzI/qDLZcOK5yjIO/Tl5TX/prAr67SS/CDbTqA4h
PtFc1B7Sv2qo+cDiYmyMR9wriH9QLb8F8mTlOCSGTeNUEu3bMqSbni8Eh0RvKXjE
VhC1VtLwz+WoFRh4JQJJcBx2JW5zXWhSMRQOxF8EgYZ5f+DQMc/z0DESDm9LD3mD
ldBJu1yR0qbxrJxxIrdf4qlS9FSWT3wMKt5b015lYwIA259aT9IuenR5qZZn0zYy
G0v8WTC1tV8nkWk3QL5gJa+pEZkOgAVru8COBYQBry+cHFrXo8BX4j6WqwYAziGF
6M/ryJ+gfW3gNuKA55TVW15rBIeJuQQktWywmCneH1uY0jDLf9ZXNHcjpFnwxH4c
/NVOluJ9aNImgv5zEv7fDrMPH4k2XuEbdIB11eWNt+g1lK/n7hQWnDtcpKLG13V/
8+dNZikncoRZU2RNb9CCGwNSbai7vRTRdiv16AyzgLhsgsZeNYIHGK0WOay++Sec
cHMPCD6KeGDjtmh9XjvaoEyuY0Fkjwjxl8yEygZ2ONVt72oAVSGiLjkujyZsnUzJ
AvL7GQIUcv2VggaDRr6znxg34RIWSsy/VmfLgSvCSuyPGpJlPrzxLRouitw2m7Ij
OldRGQih6bhPhRfSNkc12pJQx0vvoWUeN0buq454/FGCavxSDNwOQntH9fRGoTLB
MyZYOfoJheB3FKBT/L4JpJ1Z+T6R5jGuuAEHfqqXUdSIdlqXNDbRTmnRgfmOAOGH
gi1zVUq0MBl751WC+z3K4c0+dKgOecJTeTV3qwogkf5KmvgMk/v1iS2O2HaT1BZg
xP+FoqLRlMTVfT/ivGUF6gvM2X79Ok/AXBwdhBAnWFlaFwhAY06bsRUcG9tdHNkM
l8PsZp/P3UQ4XIzVKlwe7Jt0+97lhDaxspot9oc1XDY9z+GyFYGWa+Sc2RG6XVXe
sHq8E4UUTMldtw2gtavSImQbDfDD73qSFRFrVN9QBr6yJF2w43oXnw3kMuRchrG1
BskFQN7LkmzPzkxQ00oy02mMbSticshpRzbLRrEsV/SWO+B9LMT5Ovrvxg14EILJ
Cxs+v7PgbPgEkX5ARaZIblcaXJ9jOE86k+21/RCJfC5oa79KBufRvl9QtbjL+9MC
7F7ZAsTFOyByGFpaf8soOgGL5mcdrdZpztCwNNMlfDexI3G4E7VJNpGTArxLBseu
bPGnsbeESyreSVWPxADDQo/y5SNbHKNPP1hgA6WVedangconZTS8+P/R/LmhZ3CT
YlQQXjU6yWBmeOu0hSLS0SgmrA0de0BFLFvP66Wi6oq4bDzxEH1p65Cq/YOkfOOo
0ZGgWQFUfv+1gtzJhtnEDJwWH1ndzbBDPne5T4tLfuohEihX/Q65gCk7sNXjHXAh
BDi6jJYn0HhWqtQQeS0zJe7xV8ReO2g/Rkte8+f8XvZisD98KUAWKNQU8CyhAINo
UQdO1LiP8wrACY3zBDwukKMuM2Rq50RsoVLxhPCnL/kN9AuKLWeMYSK83eKPFjNy
2KYdQLr9DYEEIAv2UC/psWxBFyBl7/qbuGl1uxZ7HzMQOn2pzoYhNQwB4WSIc/xg
lZQWHIIoc2TzQDhmSB61KGHMDAjJvxXLfCrtsuGyPm9/U2vPFTaEELN674gHgZLW
WeRlRXhTGZnQkkC4dWGmH+OXBQM+no428ihJf43pyBoOCJ5dvEsv1HwlqfNlf1sb
pp8cqSILvdcYYCbIvribw9gRUMheEeRfCKjPfEC35evvTRefNr6C278n9RW3f4VW
Q4hpIdXsMV4vj8zMg6xDaeSWNZvlth4R4xQyrs0vK2Te1fYVvly+lwnPmx0ypye/
S/2iQrSr+p8e1sfkec28bv62bkE0yigCDbS9SOJnx4wVNpxDVWAuZG8mDdkVoPB1
8pDB1JEX8cKbR3nRcopJyQvAnOm87H7n/gt1s1E9rbsyE6+lZTgoXRCk4RU/Po/g
kGV3vDu18PwIu+t6/WjxeP9M3ROm66p1DLfFVVW6WMDZPWlI9gReujQWxNTTKJJS
fL1wIXCtyq1pnLSrqwj+XnVyxm3WM5YE0Che+OuKLP1/SB8y7v1V8TeSoaWZG5z8
aPPbEha/1LioybTykqnxg+jlpu+7lUfcx6RKh6+WTZhnMYxZSTri97LLTYZxSqyJ
Tqw+IFhz4IPMa74+w3U58Jf2DC/k16CXe0BVDyPKiR8aR2xs3qsn26UDxjYR8LCz
an7Py5f0PLLGSdSI2qsSANm9lW9X0DK4vsVKW0fCSo+WUgoW8/EjyI83mQZJmiU8
daefppx3Sb6O44FDJtSCZYnqL+i3HDwCw4FD9vI7/7GPAJbeqADg6GthKINnof5C
HwO/lrhxsWUWatBupjZP8E5G+FecyetzX5dpv6LbICDSex+q2FXqESDCkylAF/Uy
LEbVoahEdvTmSSUsb1hkDeDtXC6IPGFVPpcO8A/9dbFfJHZUB2zep4SCL8AzxR0s
ZTA2qdWnIomheB9fmTbNk4mxvpMtT4+0u2CBAhRw/r0Cx4wQzRrkhChzZ1bq77LX
JaiKaPVTwOv+19FqWoOOzj3K8ZECzGfmG2yqXEKWsW9iJYM1OwRhEpFayllD/8gD
0IGTTFqgj+dzmuZVvuMsQQttLnKbfEmvM4IIG8YJbTHWJZxcs/PyObXCR3HZHBB0
vaR2Eq7mAjxTfHrLNGKdQmXG9LSgx2d+kEEILizSqjQJciGnWiUhPfnWmcvHFsF6
L64TJweIdWlwW71wiayxAEmiu7VJszQkwz7ms1egC14+A2c84uqydn8jHI2pYm6w
+5Uc1oM2sAKI7XcCEhOEEItbQvGLPc4e+vFEDehJ7r6j0UtGlp9JOlcGBhRiCYo3
euBy3BOVXNYYTcuk5o3o27LhGFxrcuLD1vWHI1JyWbtoxankmJSQcTzgnFTLjwPW
aoiHDmWcndglxNrhXT7ij0XroJN9stTA3f0NkRJt0pwPgdlDRA7BGjeGpeZ/nmVR
TESkQLySt1YPITAaaWqQ/0nrpY7Opp7Lly2CaeKWnyGupm2kdC+A/mtYQS6MKEkY
AI+ewDgsrQA//1JfYqt3cIaO2sraBt8d+FhHJg/+qNcJ9eYit//jwBBTtgSjZSjj
SD0LqbTYyeWC4t+fTghmimlGnxi1uHiQxyzgRTdLTm9l/HIQxx+gk9qp8Le8Xl/y
2GzU5IomTtn/jDjRVM1HnFa08+9kBsnW/YPRY5P5YwA8XMZA34awCk8APtE0k6Dw
Qqgo1JSnHLXL/oMjlssAAtOjS7Dg3lDCe7YoXkHgI1EqnOaDqMzepDSINUh5PFT1
35dds7hGKSdA3uP1W6llba0zvzwpLWQ0ZeS3/YDFaA6Ey/BP0FFeQ6fCKdd6z/07
BVeloIv6pEkHdr7qeiPDBBFZiSrrNrFTDD19NTvPliKcjAL3SJRPRkDOmXX0OcFc
iDYImkr3lFabf4nRmqcuScooscjKOvGifWVNzVD/ssQDfe13oYU5Hbaa8V1BBtJF
a87k4Qd6gQdSCBUxKqDjJTqU3cSTP5VVVibwO9EmGGfQCTarz/9k6OfIqxJ+XON1
z3qQxRCHGX8OqyB72nCC/nD/P3YdYS3qkrU51e/owO2kvdLN+9YHC+oGJHQIcZL1
CceThHZKJDriZoA3of3r46X/ECKAaHhxwtSytS68ZL5Q53OHVD0ASHAhCb9ORHPn
0i/tkoKm7PXtg+stuRiFaoqbHna5SN7bdi9zvh8AVs8Xh5pw9sI2Sn//Bw9WZB7c
xfwpiW2GR58oPZJJG3U/TD4w74Df33QOJt/krG9tJgLHjJLXlozWAD0i67QFfKqZ
ZNI29j6X8/ZivWQPr3fGQVLSdqOSUjJDgcfSlflxaUsQyK/bDPvs79K0jbP774uG
TXT+wqUMYiaiW2ZpFD93d+sfVo5yYXO62/pULrliUnCyArJTqz4jKGi/cZN4/Ifv
KOtn20/vvOCQpPgRM5rRVwnCS7msQ52IgtWkwFSBy9VuewgSY/XNSsdN4BPvK4tG
FAifr4riXGzM0UOUZKyEtPf3/1+Y3Xjv9mCTzcfqvF2oVUc92FWhngAjnYX+dmSZ
cIWkADjsMT2HZ1ahGSAtiPkwnkTRHjKpQkxEe9LiXFi0ucGh6MYSOuP8LGbn9k72
nQIw5Qc3QZ795EJNmJQsx4j7hdFCahCFoszjaoTyUyUG09S+I/0RC1J4WEdo3vx9
aG0Gn0LeWWBZQzsiIuoYlbjS6sSVyZty31m+fO9X3irO0i4SqBFRPmQO9bQ/LMEk
2y3WHCOaU5JRWGstX2/oLg87jtx7jWw+uThuIE5h/bqKjTknDktFVcHZEGuLU4pZ
193IQLpbOhyupp5Nf0Q7drFKDUEzs0Os0Ts5leGFOfrTEmbUEd9i0l++u51X1zps
zK9h0c5uicBWu5yLaQfqg5UUKTx2LlyC/2q0eZraKhHxFKQFZeBnS5zyQJB3WJPm
lKUbUc5/sgKTKsSz7gwS9RfYWgYWvkrQEPYJY3H9ijrClJI+hVi0QadRJtExe/eA
LfCLvMUu+xZ263AWaWy4tJGgmoU4C6Kx270wON0/8YtlvBn+sVqWGKwplUY/x/wc
HuapUuOC4t5+msbmML26aJ2vVuziaJO/rT5l9COpdYl5c4l6lWLc5gf5asMQDIl8
utyCUXKtzA6D2bS5FtGKfstgo+YeqFTZfp+azH2wGFAK0/81uEhEiPaKS82xG8fh
zzIGbQvQfBFGE1I+v8LTLx0Jn/pPmScachg1BdfX9jcVO4RSLzZZhZZ+o8T8w9kd
ysmkYgQb0+acOIlKw/RyCyw86xPCpaCv1f4k1u+T+pQEA4QYV7ClGsdAzHu/FvAG
ipWQNLY5IR0YWkQjUFDFpkLWA7TeKQov5LHVI9KTpfkDER5ofR1ed5LWaTgwkPU3
PJVM81mmXXcZtMeZW1N/BwUWjL7DL34t310vlf4iVxkqAAVgUA9kJSySq90pcPWM
w9VLyMijc4s//1k8a1ymjIlC7oJy2/8sgllyZJmHJG8Zp9bu3am7TaVDOdfH0hMb
PhYYs7Wj/NCGy3uHOR+zQrRr1Su8atouczTL6ShcO0Jxgy0NL0yKD3fbTp8sps30
Lc8CD8IaLHkSwmu2Nk+BGSMmlSzNeJ+GXCpRGz4jpAb/6MipmCuJzEqApFp3Gk39
KVgygbB2UTUgfNcjk1BgZx+TsdL2nM3tMVqdnHoJga1zQBbXKeu1SMWqsPkY2mSg
Uu9edgJmO62ZbwiFmC1sKasz54WD5Wm60+KX4rc3+9S5eruwo9kZEAra4EDPE5j6
Vq6Db39jiSMBRT7iIbVuVQfAwGbDQkrGM+YeBoOwA0efpfnS0Cdk8oUjNhZ/0NSf
sxohVmNUcQgQMhvquYy1G1rN7EpfiJdMTwn0mdH6e9TxhhAr15jbryw7GjonCGNl
hTh/GBbWk+TSP5d/x2KsfNUPs82gjZSSqnZAtbgGasR6FwwLErZHuF46a50cqi0w
nnTQadhf6B7oQbh7nkfIF6LvBRYxuSZ5ZxADKiptUKZ7Fm9jrGzvcAS2FaeTObol
rS9aTB3DZh/WyWublvmx2K6e8KBAS24mIVKCbZQsFlvRVzNQ3W4092l1NQOdIYKi
VnjNdwqPODDcCA/b6iozUcOmoXcahReWXTlaL/KE7csxacgKeGnbrfoMKhpnHMx4
XAVG3icmFFmOcMhMfpZ/6JpmZiu3vrPzgl9UdaKuVGYJiskDdmDAslv3GGKst4B+
fraWaP7wHQALcD6RFK2EMWMR/kc36lZ27FyOoveHBopuYdBzyjDrG+y8QkFcLqC/
8c2gFMhP2g8BxCFi3Iw8m6gc6u+nEkOciSiQ7i+mhXszpeMzEHYfc4r1waZ+K0wo
lr5CK2UQaRZwfmf/605Fhuej8zTU+9VPQ2hP1EL9YzkF+lRsYmLfnibHs0sRyYJ1
xLqgthFAc4Joa5aLnG+0KpnAJljp2puXw94Z3ULPKnmN1E5/ezmSR9ArbnM7ADhq
WiWtxuZDA38HYQc1i7xpFteeEVCvr1ecUsE7Yx8QyX1kB4i+Uftg8u42t/7DY7sh
b6aDjkQhvUprbKI2rAjjcwIJTfBZJFV2MbXW0WNmQn6q0glfkAcfXLzoB9UVLooP
Q6wKRD9yVYlvXny9Q8X+/u+J7mnFnJMnwcIO3+/hy0MEbX/BmW1sQwn7ZyFOD1yn
nG7olns8mbBl11xV1ocgUOkUJ9hh3VtjOys9JtrMU3Hoz4XB6vsVgxKkhjU1J2+W
s6lT5Z+bywUniVAo7czmH1r4o7qFvHOQlUOsLU7tBq5B5kDq9cSwSWh9HsbVdJUd
8yatJeVX23CV3E/3PdI29eYAf0zKLux5lgVtkvcZOh/JEZGb2F8vU+ZTwsfuQae2
U9TDz+uoJ3FsJ35NRkVHN7VbUbdDkAM1dhrCYsHaf5bbmqVyh0x1HygYXH1F6Omo
XeBdvRn7bkFHRwnYLS2iQ1S/Bp4O4At4g0eYKn5Ux4MBvMlw+g/SlgX+1SHSwSyq
YBJMj4nryCrgzm8ZgGW/Ud7IdkzYBck9eBN07y0zLx7K2ResSUuoGXL1N4iARTqn
IHyBkR5xaJo9VrOeYXmO/iC53UrMN4KJntsplDaDYbyTMGBECc0UFQnoBh/5LVx8
Mqgqq4l0YGCwp6I0agaFDybNjC/NtGB1xIubAOLjjSZxsQdPBueVaw2ZvaaYLcTT
VWmO3clbd3P9Ief2CjEDZKZoxW9N7BYRIi/6vWa+oNfhzM7IzeWq+D1062qrFNt7
95n4pOj8/TqTXm8elrBQGrJNRMxy7BW8F8RRRJmwQYVBgs00cEUworBVml9lVsGI
wIPyLNusN6GxSaj5ZvIg8VFxDY0rxkdyMVK3AHwhjQtLa1qpvRSUvENRf9DrHBt0
qh0cB+qyUIwHoEr8CJJOSwIn7iIGLLtDw1PfT1STF0GntWxwysDg82SExs3owHYa
PVKWM8wPahBvDEgI+MuycSOpu4gVEnO7iwU+5YkWIXYDmcWNGEnbkXB6mByVWPv/
RU1C7b+YxMKfIuJE8o9S74AGR9A9tooIVYIayRZ5A/eknx0O47Rx/T+Gr9VfNxHD
2HhSqXzm7KQ2hzTKpEg9HHpekz9CfnPORUMLjvyC1XA0L4fxVhWS4CUN07ACnBvA
wE3GpXcS2BImpVPHu97gOS3O7MswymRRIB4UHlMGBmt0teaI9LYYtyPqc3bhUilj
v8jOvd0Uv8fy/oK8tgZtSe98vPHd2TByhxcnCb8jn3/4xat2JZnd+SKpvlA3zqc7
Ac2BiEL4bHq3UH67HNrAswOZ/Fq/CHjkrgRO3kQa84VuZXdafiZ+EOKQ6MHu6fR0
ASWZfG7ZX7JQVYGyRUCA9xyMxTKOLBmQRn9+jryFkMgXK9gPAe1TrmxjbLKbIVIQ
Ak7nQMRJLyIcZxF8MbFXDLXGzCSAS8P2cYNHB+msxEbv3r/T3tPeq/QEEx7mnkPI
hS/hosxqG9Y8KlDimGZa7l4PfEc819KB6wMYrttAn7QXfMZm2HuIqdlEVVCOymfQ
OophSgcBUwGnypvlkje1jLpfCkmBCftChS36Y02el1q/DcNvml4jgoIs2yNvDCNb
PzTQpA52MnB/iC+90JR3wkS9Y7hh+WH/lZVgRISbvOG8M2QNK+wJwOIXMGe3h7Sw
e6Srb0eow+So5hNQn6/lM8gkzqmwKRblMVYDwbJhF0V5E5Sqkr259mf+knsHSxZp
Zx9qXsjFKX/V3gcNcJ18XFrdpx2rrL9AFvB+Z8qtFiAo/zz+LH7oyqt6mz2MrfzB
WVgzQrFwF8YeMp9I10ZO16cbVJqEwOZ9odcJM2UT37cUiAN0Has5ApXn31v5EKex
3jDu7Tr/+Bg4xg+0w3TQC05pLt7X8dp0J7sRMVqw0IWfoSm+0l7ZFTaKEGgCJEWE
EKqVVzWSL7JE9AUdkgIsi4Ta+9Oq1rg8A1jyhjcPIM8ARvOrxBfq7ARI03jiww2s
NCkrkuJmLIr20V9SjmCGH8UyIoZKlCCBaDDbe7ruQAvsYQD91AkI4fF8hdSDvuhA
TZOg0XrQFX7HTgKvKzgWfcrzLquskc6C/cVPNxzLBRUI19RcFtOiaEeJenXfSGGP
XWLA/f/vwbkmEoZrQ0JzBvd26TAZjeEusV3AKCeOa5xFoBqXx9+FYIBt3Z+avm5T
4/kdggwqjaSeqynhK8B0JMv1cwfVvIVW36RPmYNvs/k9LrDUdi+zfr9J5T+8zPk+
spYfzQFHZvy8FmKOgKJAU+RiGhU69bJbYC6nY1hkFZkD+Jt5MkTBs+9tF33N32HO
wmFiIPOOJhUnp348Jk0WcfgBsW9OE3WT6d7LhQ81982oNPdlwzvvd8AYg4tAz7+q
c9DQ5wJQf1Sdqs8fogWF2Uf8947/hpaDSrKZrtkoRDYGv5uGZodmJP2YA3azlgFe
cDU/R0r7mDEUBKODdhv5om9LG7An/lkKdk7+3qvGrUnoIUqcQTw/lGQkyvS45cqc
PLyhzVpegRcHIisx384audwd3xEUGHK8yuo5ZcE5Oa5ucpGWAmooVujXLbGPKVWZ
PrZpxGWtKxn4GthG4UKpryMKYWEeOg43pzKZFC27BwTVp58PsFzDn3rWRFOJn0sl
HIBKF15t9g46jbZzvZY1h50LWVbLhHbGKqOZzrgxSj6H2h+KVwEt+mjHg8hTXlb5
OzOJa4SIiCflR2yfFyxYViR2zB5efn4/HlmFIWlBz6fdFDIpMMC3bjzNYQUy3dbQ
YPFfaZ6Zc3C1Bf1USNdl/oxI8N/s8kpftE/OxceAKjeF5hoC+eERRPH59MhD9I0z
JIharZcKqmEyuP0+lVaIY0i2UfTqQQJ7+I+fkh+E4RNTKw79gEeZ4+0Q/Goc6eq4
Or4GZxBSKNpxyZHxw49uwFkVKJiTMf9T083pQKbBPzZ0nYi2HEtjSxuNK82Evlr4
UOoqaVVL5Wi49DyxzkiiJqupdZBybIHHo8Qq/Ng+2pU1EVfQugirLV15V/HJxcyO
5ZpEWankdfo6WO7itYx2X170BQD1+kJY8wxj6otVPQjahEZQt4i8KEkDgwF/p0H4
B27MP2UhNVcrZ8zuM4POXcV+mkFOb3ZdIe0Usm9x9rvPbbHbPtSLdBOkZ7Zh3TEB
Zkc9SuWkPUKj6HwcoLOROqJYt54zHY7kM7tqbRbiUD99tgd3qwoJBQJTTKIy6/Mg
UZGT6DF5QXX3NMUEmLE74AxRxvfbXfEmVh/nZse3g92f/f8Xd2Ww1G9QiXNd87MI
Qs/pZ5XJH8XxPE+ZvKze2+USeUsTVPGZQcx/5VHBCBo8sqrHCeYO/0K2GWouTbFf
fBC30hqRfyiUgj3vkgQBltg7hfN71n1SQFYemRmMTXZuha3Jj32As0E/MRVMShqS
7u/jNgI6jyO9P/e4ORpMGx4jmCAxd3k8oEvFoRXwbsH3B5nik7l6sOJyOj17dbsX
CA8Bp1qhyCIPPeApEe5lh+oqJZMIiEWweM5F4G2pl220YiJn5srtX9qJS539bK/G
SL+Ks0qoF879nOTd3YnYGTp543EPe3enxwC7nAkPN7wjfRvlNWrCbSpTXZvXKj7t
7NoozwV/MYa6q+H7W6ws1l9WHopkwd//7Z8GXxVbeLbgGtvuXYtBWCw1kE6/CBfg
T/rg3m9zklXVdAFKCstnj/6odzk5Q/xrO3+A+jtuF+kR87ezO4BJVq1WfVYadyd5
vEh4QLMCAmm8EJ15EA07i5afWBtzwEWp8i+BRpFppM47BEnN6Ws8zRRv47W8DRKG
ovLylGq3y35PmfzKlzCgfNJAhMRGSDcqruvdr6LH1lbrTj2+djtTfMAp2PeAd7SD
ixUxbyg36cOfKct7sQxE6CN4BNr5Q1xI+0YPequuC2JTg4LJp20qBKgTxrd/Qz7N
E/5znE5RsVuNZAYa9XEY3DyUmwXw4lhJZnNa6QFgT85YGh8wZoAL86PGtOiYrhly
NK6j1A8gG+09azKJCJW5yQdMTrQ8p7HndyHDRtWetCSDWOCFGaiSpaBR/c+hofX5
QmN91Ti1RiZVhs8aN6ffDgOhNhdYpio1vEIgco7qceHqLjKIyZkoAMc3kxTX77js
gZHlauA73tJHgM4VXIdbnRgriJznTrXtWs0JvtKj+mYlASm6PkaEwcW9ZQ+ohPJ9
PAfgVHIJLUrZuCC11EaRU8vAq8HJ/W98m7/a4VmHKfuuqdO2P5zMQGLUnySF+NRn
yZ3c+DmG6yI+6nGoBGvsYRGmukk68WY0Zx7zI9ddw3GMXb+XW+joHexIH4D3a2Cz
vV/hBdQ+DNj4tdMxvoRXCrGU+vtewPuQF3J3EXWmRlG0MkLt1piy2fNGodmliWnp
+dHiy/ePj8A5T9SuZumHemHYI9MuIHQGJqc/FzofMDPHen/SLeKUM0qu3gjLzkxi
wFZgwLsbVAu3pDqTlI5oo46Dvcs5aZXyFaU2nSCOm0FOcwi1qpUjr8pN+qEkm3gd
v3Z8plDADb4BMD9+2dD7cPRhkV04fzNf8wDTHGw/ZseqbuLsBe1iOZBIe3olQYf3
brC6KzCqzZiuZeoBTUJB1EDAj/PLGPx8QcEYa6hd07zTrHO23Fel+btwLqvY0j1x
1qX88ikeL9uOvFM7SnKjI3tj2f/nyKjLmC3jdEOxk0WSskIiM0yJM3LAJgFpoO81
bQZ8dGoVsqvbYT0YHWSMrpsNMlqDXbw0uaYGFqFiZrbvxMuaLB7L6J8ZnJvxzB/X
ZA9/oOoysDv5IjcSLRFoO+EtrA4vlOVPRxTpNrKXfrBbeTTUYIXvCmA+w6zetAVi
Sr6igbue9tExx57UkQQHbahdQ/FFqEGZDzfnWGi2D0nbKQmR6Fs1BIiO/zMUgktd
RzHQeX2+krt4OGEuWEASfbNtR+uWPw4RXq/ZFj/jrmLNK87kWR0B+arjERHJejSI
pb902btWhOY3HfDSA1U4vP7uqSVq/U2dbXp94pgK48EjRsPfuPkyuIzgU2rySYBZ
7G42F6H+LC7Pz1bHZ8vjau8jHxzeyrttXHXky/WLOTi/J+Ac8dkAGO5K2KJzgiu/
e3QqJVQ5jbBM1kIz56s6B3JiMziDHmjx+8Wi1xt7Cc/xVRDCQb9/Dka5mm2KyOuQ
m0W3250DqwDWLwREmGFfZQ0tckihLNzJ+U8+v7UfdQ4olCtwXfxvLIeWUwWIRo1E
yXYVtSRcvnAymDeSfN+NU8Z07u1OJOFMMyNRPsuIupq4l4UhVGZy3q8fnSFkAomv
SpVBB20N4/R06c/N4kAc+ATq85mIXOXFdUY6dPxQaJIvKYBp9e9S0hWIP303qBrA
wrFbqEtzzcC3cHILMWiI1vLmfQ3P6WZdY9xP7kVAAgISZU52LAjQ9cOTo/tkOKDM
zKWG8BKC9mXueVf4ipD/rbdwDzjnqlHBF0AdnRF1DJWXCB3dljPbmPHU+blr4xqP
Eldan6T4uJUsEOQcmMWUoC7RXAIQX3aTpuwcdJThkhFgonss2gmd8mUgauqPNi1I
xHQVFw2Nyn2IbzqM096xzk9AwTk809OnS+mzFdroEfe565CqBw+tTwsgzKMYIYXd
mRyVIXD9T8r5Y5vqTY1LoG+BMtKRV2OciZ/sT4iXUHmNeDL7Iz4jRS47TpmdqotR
jcyNMMw2KU7YTIWUu0PEurDTNVSVsP3S+a37ghZUrjjsc4WceVXi9sT58LzEuj/2
EbGX+UrDrHwvZ8Ii5gZkICJbkxmh+kUhFVbO0y9DWrgv/iPvb/n9qxUQMZbgiGpy
Dzoq+SSGOCdvX3IMG9n9jpF1WeWuHsH43xs4BD9/s5vZ7qyDh92DT3QtavRpKu8Z
rEFnDTDnm+zQmSWV+vXYVVMpSV/tE6v8syLZX19OXQYLnm+mQLV5ZOA9/BA7w3Ke
r3kFwCwrFFcg0ZYPI4zTP0spT2j9rvYNRE2Btg6Bnllkc3hJEwzi40tPOC29vu/1
Mdy6iOd2SlY/Y6KUIq1iHI/6G0Pg5dVHb/nhcNrQCRlrFNvDOw+MXvFWaR2JA6Xz
O5/fxL4cATnkH4TcjxUDaCOBly6fZ2j4bZTw8/q4UGsaKt1OMRTqQbrJ1p8v/UY6
d7irNE0xKhDpcsvKGaEdQrYBHP1zTlI3I+4QvNdumxV7LxbE2uwJP+XHxpqwQZVk
gIIkEfpai7MqDgPp8aNLJlHeqyQFJ2QWBSZAeNMCKQ6yCWAE3ee3lMp2nTzMv6Qz
nyrUl39vwavW7DUgD3omHTtg6WDhj8kl6eEwiB4qH+6lrJFbn8spYrnJk/0z+hui
UtcKLR5l8UUJumGlLTq+G5uB+CnpPlRhZpdjdFsaggncyvQjUomQ2QP30rntIVtf
1oHW19ehgyoBVFp3yVwpMvj3pGtpQ29nPnbVuFPAwYq9HVTWwNlNvRXBXNT5eiBW
JsJNSxrDSO+j1Rsv1zkYVFBDvX1p/4w5523xPmjwA5fanCtvrCiIbMEQIVWxhR8p
EuUUUkbAaXRzWbTdI9kXOAWAR4RoJcig9qDplnKv9GhGpGWF25yZ/SPxq2U3pYpc
Lm4YBT08BYfcX9y6GoPnQzz++IwxKstCphk7uDvxn84fBiwOeZUyT/ZUvlE6PVSX
FqrZPp4m8o1M1NMvDi9O91fswEj1iGcopGCGcz2jfeLlUZro37MOZGjgE5wtn7L/
ZnsWg+n+znTlJV4v5wAGPT4093snj6bO7ZiSx3KoQd/kYPCkyNTK5r6A6HPTEJQJ
T13WeNwP6EVwneM7mqC2bhyT1u9H9Fs+pzwAcMepAH8r2lodN7UCJvTzaOUHdAxp
fDsdm92Jyd2wbTMGU99soR9mAk5TUxiBpjmG1E81EWOcurNcD0Y3Qa2ueNU40Lhs
r/O3doeZvOYNUoBnTOd1pesc7Yso0+zvJbmtMb9jxBfvNPzyAD7hv8xxae55BP8C
b3EsZc4NfkTUrRwV0seYpXX1CNNkV/VJvSykZ/+5GbfYJ2eeahqoPj5ENLHlW7Ok
2+LRCJmWDEo7aN9uc40flYvcvY3Bo/vSwIIRbGYklSkJlnkh9/RUZxSohsGflahf
gS+gMmXc1ZcY/j9gwIBOHXSpQTvAb/uR0zM8tCafDCL8cibNZbrWwL3E7/7pcFoX
FbGG8Hg92tHzHOrJDrav2Z6DkKBwnX4IoviSG/gbzS7XSlvjNduOOjTTb0Cstmnd
nbRlw0eAouVjPD+LxqlM2SuKea0F+Z/9NiqrvxaB+Z96kYHJQzEbwu94wJG/wUX8
rGSTwQSnC0x4NCeZxFC71/psY0bPMpVCs0JuZU7PJZnnsH/mt+TgFHWOyZLJAJ5p
Z1QFmlBm/fQXfL0Hij/Ex3IraGNeIQaQRZRKqPn6HUkUwC8cF3mjQO5eha/TQQeR
AZ/2t9RZdWK98v3em0cDYJvo66VxTsDw8WWiyITF55HN+PE8Yx1Bin7WGcLy+GXj
vTpo0PjoKs70TeQ/2NBjzQXYLLD0cNmB0eRSBVsZSPwmuyAq1G7EAgdSLWuB/CU1
1rF6GjRwBTFbMdwG2xlaOu7SjY0StOnTgxcliN9kEGuWXlX3yjsI1i4FWcMhLdf+
B8W8zc8yg9HjFETWZ4O1EpC0iTFi44G7z7Bvz2i+AfSvou42bNYCehRqUQtG/6FB
eGynUzPFVXWZuuH9SWbFRAIOUy5F0nXW4zxQfRHU3/fapHIGN405n7thjHPMzVbP
jgSYoZHhVAUnf2S2kix1E5sM9BERfcuufawRDWQ81hEw8EH8xG+LRibdKNgc8b6x
wC5V6FFZW10nNjbS2z7ghoPp5jJCud92WloxyF02u98B0vg1WB3QIwS+I6ztX69G
L9WbksjExn4/pLq/8Gf1GdZH0UUX+beaMTxY7GSaWFQkG5rFabbeS10G92W4X2QA
2jG6sx/kR5dqzBHsS7T6YjrXqoZfYFGD7elbyG7OJFJ27AcD75jEl9RyZDGahB2U
zo66DPF7jgO1vfj9sgANdf7dF2n6VRKTxizCmqH8VCM3gE/J4Z4c/YB+qV+q3Co9
7nfGeQbmBgfHOwblKlHj+y9hCfJAbaJarEeWtbXLzAsA+iuozBeLh0FPy56SlsP8
CBjK6vyhYDSZ4gobeKLaEg8aQ5AB6QijnpOU88xf3RxNnw0xi63ng1pSJxaByfrf
0ftcdK+M+PWwJhwOMKe3dJtHzSabR+ncvG+GCuJ2WJWE8j7V1Q6WtJqWLvAyxfVU
dMluvl/vhuFEP0fi9pLnZpG9xeXlN9k7DNdL/wRCFPDRrScjglwEmO/99Q0MiyXK
ns6GPY06/4E44z3nONlNxJ8rxkt/t7/+di9n3T9Qy4kB8/B00UnDv4PysL/3DoKf
0m06BjVje6zGk8tjDSRasq6gjHIna0gBrtCGDd27OGujt8ztRRNCwiTahbJhtfZp
PbobwYCfEEY+LieFGeHpDTh10LccrMSM+jIDIaq2MAc76G1vicu+MhVjKX2K+4BI
Yw/Mp1vORRc98nwDsWg8rjAOn7yaWku6hLOWSmEoCdaQ2mn+Vh19bxrJUD6w9Qn7
RYtaMgYNZw5ZPkDmRo/6od1SNbarJ7qGOHBE+Yoi11hVxfGFmx+JxxQ4U7g9+PpO
s4dlXaSd9xCawEEIwNFQxFtRHxFKCOtrEED4HoFHkBkW/332J9j1Wc7Kd4Ic+uyo
xbOg/H8ZEdcJBmWOBAYQ/94qyqf4D8a+4jc/XxKnMsPhXFKXVL1PWvXJO9JuR+/Q
9JORwrmYjgjbgIQI3bl+XTdN7XzicKpAqYeU7ym3toyT84CuDrrmRTylorbb875T
8pDXS8KZmsmpW9pglffyc22CnVN5dLQ/uu9BLROk3owaTIgPk3C651DYs9wlWH5Q
Mtviv6ldN5VNs/n9/ONr6sigBWCUY0iSfhFlVosLk6s9uSJuQsTEhgF/PyLg5U2V
lDZHTLWLoJfNFC3ntvsIk0sV4sLPKPus39vLr/e2nrXkpmV+wK6/w7mnur83T34j
LWKCt6gNoxr8Mv5aZbbkxxKcjgMjEnWn6zS5IuRKMztUwAfWWU7lbZofMWHfPmRe
xbjf4uPmB6VbSq3jYj0cCX5CCIimyj+qT9WPtFGcVx3K8ZwUVaYL/Eer/Q6IvmdD
9upMrggzYq9ZM4UCgfUxYqtAg/GmeIgqWonvAMnlPFIG2+MG1epQeq1jVNhLtkkC
ZT6/w1KitlGngNIzptFylgpwjXuAe7XK909ESkAbXtdoKXk99xtc/bsvIDRWN+NV
cBiBdJ1W7VQ6tCVy5H7C2zJIk6xjh0kRKq7wOm9w1Vm7GxMGHaYcl8iZMnu1Bvcu
g85mqt/EBHmR5lm1pG24CmOn6KQm1KKDAIZgcIZZSXCAx7xK1Zj7eJfzKYZlOZ3u
ADoD+Xdz2NkRf6eTr/4aDNtkI7NIe3/UY1FAC0kF8VpDf6hsurANT96AlArhJJH/
hg4TqolPqdcC9VDtCMlGCpanuxfITa7KuLeVL3zOu4XMwVnnpt5t2jfgFf6K84A4
iPUvZpde/yLmiQECvdW9vquGuKbzrCKCadPrNKIqLpKcL4LaK63JeN7eb5ksyuzM
JeYum+9yJWao9MTzrXoxAj1xk9HoZdLbM/SpR2bj3j4STzgueIw7VGYb+kIkQNjN
HLO1P7K5AVHXQRJ14NXboQgRWp9d5mBcD58JsAnFF9ap5KyOOZCuk7ONJ2ODwoTn
wht8injDOxSyEwkjSy3Ij+5awaTEvfHNlWZd729U720VS6lhWi4yWC3HvV6vmN2I
POP2/Y1ZqdYwBYV+vkVH5UjPsfNZpc7T+AILUJOy2mvAKf/LXCqXsnArkbsbpKno
cfgAP5PP3JvDFTQ9AQ/rTPz7vw5Onj7ZJaQ6qZ0B4N4b93fqTclhsuRRT3u0BDsq
jg+pIXs+RY5ykNByhifF1b1//Gx8k4NlAAQ0jRZuuLkq16QoybzSs7E1/6QCuxfi
xT4+rfyFNgJI+62hwS25iwytB3UAiNNuHgfu+ZXBin2SANJgkrhHGRx8nUVfJo0T
JRfc1jQ+PbTV8AfmvOT35Dh3V2+JZ/xt6Los+o51rB9xODsdGoJdXv1xdhrMgqbR
3xHJjUr11g7s7a7IL0wVhc/5AqtcaNmQgpanw3IDd3UP8K/10FKx9bvzpYBtr1On
UWb3zGpeIQDsu6jYXsOwuxXMA3i/5wLOtmk3L5hPD+nPdp85sx0e5Y+sOUyNPbGT
9Ri9fCF7RIuAUPZN8pHxLOZ9Mu66nGI3gKKcsX4Y0+Od10LBLQ6SLJvWBotSrOMa
qYG60NZTC1EjR1KGWF0kAyH6/tFlCBrHKWvQM3l9xEyYNWCC5DPz4Z2UPVMyRQYf
s5nhrNgwpz9hCi0yzZaZtLuTREv3lL2DO6ZneCYsqlB5aU6KOwvr+6oiVtB8RqAi
cja2GEUCZu5fi1x0zX2FdRMJT6cVoP1C1lotogw0O/z8Ku92rnIt8to7Ly7xCNu9
oAc7FPaCzou4FpKSxYucZ8Q4sssjrr+cjWdRuRvijjfV4XQA1bOv0JuDIWmizWFD
qKSQ+d5t0Jji0lHLqnUDAQo+45y1czKpjvSNK3NhVcd4pJuvNKxaXb05sKurJ/yk
XqMi5CMQ/Kv6vMDwzt+rH6MVhZHb61egYrnrwVEhXubAE8USiVH5QhvqPg85fbV0
p56AL11LMbZl1rHUqhObL2fZ+Xp+Y6pY3LPyxqcYci3M//qfKj+wWFDCXAhUSxXb
+DyqScc/LIBGmLq46zxlwisGk1iX2Z/PhIAFwHor2E548zo9M4MAVgshhhMIUi96
48QyvWOsjCcEFNJCq/15mzPS+Cee+sIlH7ejZIrQ/fCxr1KSSkccx76DPRlQyI2o
tZQ6lKSwAMuLD+n0sy0MnNY06OAqpuOsDChto8weUOwG8Nzlm3ib2bHx4AS6hN+R
lJo3+QcKiLO2xlCARyI4/2MhU2v9ainfjaugsij8SygFuPQMC2mEmiTCU/c9hATz
P2x/xNeqm3QfdwzPNHmUptUTO3PU4ILuMxDevCFIW23PwcnVvaHEsFbykCGJa/UT
RD/R7nws0VTPwzpFc/cd5bLCzx+e9Y8D9Ur1WAzH1WaHg8cHqQmWB8+LgQUPq9Gk
iRPlI0WXrSmMj0+Rm4BBgVPTwYV4kj1d+0aHMdYMacnpozSOI3mILox9MqZj8NGs
tDKgv5mLLqkOzHBCTPw5j2q6VhE0nvmMiiC3qu2EECqV308VtT97TbFoDx3S5gwB
euIWPplugdc2n/7APUOE2kgEF1L8yXmK0yM4IjYhdRMhSlthkCinmcRxrAbbVTG6
cVp0LTR9JVAvz0ZyV87LC2sSyVShLdmajDFpT1DnuGbTbcXK4Ue4ilhKMiP+UZ65
IivsCJvi2l8bDBSPL4/CA9PK2O5UUPf3usfhL5qE84ljuDkYN3IKVXjC17io6zEI
pWovVc+C7hsEbpArqpmYiiBZl0BgA0tBiDz3Ws3X/i2qrnqc69mWrPcQum154voJ
7nDIjab0342Tr0c1rQk/+b6iU4YJBwPc05beRiyeGhTj+NbjLuQScNTrjXS0TvTC
FUvQ0JV5B8G3h88v5Tm8Avto7I6pNptd7KezDZNGagRRyAO30EUXRdYsvM9c11lm
UhoLqCf3zatZrNBwa0RRyKbLERYWsaIAo3sb4JYg1EbndJEpRvQccUU9DOkdTgD2
zeo3WK4NtLNP875WlsHg7FAYcFIFZ35RQABrGoqbJVRb+2Afz0mcgMJCPYwozbjI
5xMoaoVr5RpF9jUrxmcydbZJQskf7LSd3sts3G12RPrl9d20hpQTWegxt4gCSwxj
AQ8/Ie+h1sATi2kdAYNy5bieShqv6PN2kSOMmETgDBfaaqwBwMsykPXH5Gj00Q9J
2Ga3/pctUbDt03qWavmYsuT67uNHbGUzoPA1+zdFd0w5S+5NLgrFBvpY/JyMi/oi
BuY8XZI12MTkE9P0qpugRz0IgVoRFRtQ8G9Xd00VfSAokYl996dw87eANIizjJDt
k7O1CW55DxDyQz1rbkfjDggrtSfjtXow6MWmYhyVuPjbdbRn7Fve2WYJjWc5zepS
j8C5shBPBLZJZOV2MOoQRs0+o+WrUovNDiaQ+AK4d3ftTYzBofwb7Y3XYUe16tb6
f596IoDp4H1LtORAdj66kTt4bb0pZso3LcIz+uA8F2onYn1QJsv7idH2/RqLvOhI
j6b9ODPQknKvqYUBguOTyeWAni+/ikgV7Yg0XvKEai04olWilSCMbXW37M5rYQBL
Vs8www5Ia0sMcDWB11eGnuVndG19WDqBlDW5ZPckTqSP/8k/KzJjasycQASEK7Fe
UGsuKiJKylQY/K0DIwkBBbnr54peNONJ3O820KDpnznmPPgoHJGObCo7i6F0ipYr
3wjFe2XqW/IWp0Rl7FXGhhhGWfcwo7fWF6Xh1qLAtMCeiTGSeehNt5+fsTVQNHep
B7mWxtr/Ti8S89rV2nLGJeI8sT19y/6BFHomR2aV9y4TACcLHDVdMB6rqoHIeROo
Kvrf2cuTY3ONrVuojdXAo5lnYDOPCkYQw6DcEaQnAx0SaFUjbL+QSKxFvQGWeM5e
l3AxHCpZXQSAJEJIrmcS4//Rg2zUHRsTKEB39wMN2GTGKrK4gX5c7mOqrzFOY2qe
4gE6vUFUKFTvxi8jHbkk4ERjK2HXIjKjyHBkBOMJ2PfkYMGhXyQtYi3WlMFOHlxZ
fvZthSnHw3X3LUqN/YR0dyKLkXr7TF8gvPUmx2bjNSVIxKO4tKVnhmJpIO7UXGq3
QBiscyJHsPb3KPrgl1FhrZi9hQUnfs9nRAHvt0fTHS6cDqddLIG6U7WtupQxFy0L
rsNpCfnQVBt6/cPgMHee99ZlkSr2jqeeOko39xqdaRS3UWDgP+uFhde7UHuAqlkZ
ZWkychAb0fx5Kx8Cy4QD7H7kfJaeWzjjEGEbrc6jY903yT5YuxYxuufyl/e//FBh
4ih3AqxM3xifTZB3Bkg4upcQsFS6bTpfdRy21e+aKXhizTL4rMRVW4eLqx1+VSWT
TOjBIxb4okUadpdpkVrx8CQBkUD1aIfignGxFgfLRSdfV/H++IBUu/XhcvISGCaD
+aAWPTJ0+lgWe8oW5Uba/tJDd5kBRck3CfGXBV1EyP59XnnomW8Hr1uJszYetH+G
1xnN1beHx/qsFIj32j0rxzDC+daRTgYuDwn2S7GIzpB+9xloR1LjwcwgK2x0/V7Q
+YVoi98kBGnDTWZ78koHytBmFeJ2o79Fq/KM75CBOTmpd0Xxs4yqdYNONkn4bIRz
1o5Gpn54KRBa+XB6o74UssJBY5ffeSBBzx3pbsXLMdBBrUvH1fXP0bzdbtLP21Sd
3RwCvEmJBaszWLKtlyZhVdzjkTofH3MJupw238u0qrRIkmvcJKvNYGz6e0NyUtIo
iL7vWeK1ww5o6DLouwiBQNuH4c7GSDEgQQdfn7eHeJwmsUBfRhxpAMqDqARX322Z
dIaW05+B/imFQFseqBePjY+F50fxdo23RbcqgDffdAVY25yVOzO9RSJ9HvW5QCt8
tvGvS1KmaoEWzvvpVKc6EVg8j+KgFh2MdAdHtbvU0KEPCGOuOa6m8WcDRrvqDOMB
jnaZMSBjW/jS3UNZppf3mtNm/iHWJarV/XoKCx2oLEsibKxnUW0j0Lqa12elTSSq
miUbGMKwRIMILRZn/iekwXoA/22ROHIvd2j3hV9HUla1bW1IfDskZngheNySgbzY
+eXn5s3NJ3QLlUZgy4y/GGeNnXbPahHmLFoTu6TxOUOqAPoxlO/UDof+6XITnB5U
wUUfFwO27DicrIo/aU+Axo7Kzs5YdphjsJ8NJNE+4Vi/DO6JXee8JXNRv6Vel0Sq
Epz01Xuio1aW2QFDd8awHMPPy911C+qpo6D074mclCdbklAqbc8OuvSrr6YkjyAw
cygdYkKASrSRDLugFRKsha6TbzRzPtZ1MjxPYH6Pl9TtNjJPka0GAUkgpcZ907zm
NWJYETP3Aby1YgsZHCs2FrmL7ZhNtCLeq8wNf628OTGYKkgbcqUt/NlZLnPjyqIq
xGGoAOyNU4rrpL1wulopJrk5plScwFcVsKYJZsKJx8iXdH9T0rVPQpVcUajjqk2J
fPUlv+vEdgbS0VSpspZrjqrIwQTlrXtB8kqYM5A5RSGX0HpLoopMNm4KtcqwzVvE
/K1EFUIYzvZwzp3Z5jICcRGs8/XKnjgq/21SJ4K7RFs+Wa4qWtxmrFgCLr5Z5NCm
mXU+5UOjpPNp8y846AsSKwMo868PruK9r5JSYHrAb/I2ATWXZ6CSKL+4ej0+7xjo
igo9i3sjBZs9NifuwnPmsOqa9AFEVgfyTw/4hvNb/7KQioFTFsis7TGiXzoLXbrC
195mvu2eXEZU3cB8i7MT8MltUSmSuLyNc2oXgbh02xhRO226tsMsx7q9oq7St+cD
ND+6HAIryXBNYGqpBwTffioJK+Z6T/YZvMxVaVhwI+tVMR4QLJssso5LZ4Dr8DEA
WKrq7WuPjHie7LOvyCmnAjW7ipZbOD9YE0K3WLgx+FftjmeSpxYcbY408D+ECt8g
26jwDhf9gBjCbUN+V/nvVYu+PeaePqgCtaUm6blbSTkLrvOl6mjeunh0jDnZt/H5
u/HeToEvcUKtAbLEAWjojaSfhokFf9wL/vXVCll7y45HqJcvroxEaX5FFban7pDy
V93NbaS/QJwF4OlxmK2Z7uD0nRmIV6zh9wE97yhLGi0fMkDUdYje7caqD7TWDgoS
LkwCRBUZ5P9RB00qTnqVuYSYjbwFYkyc3S+wxdIDXTCTzkgMxY+74sMpxcDzWEzz
YT8sGmp0ztyfeSjN10tQXs7Tfsd9H1SGIe8+8ntzoGZdjKI0JMft19n/Vzlwd+9M
KBF8J4KCdEHsVZ/i98V1WsEWqViFkupFqnroeNI4gstwhvPeKQnTJnnBXdNEhmRD
CsJN2MDoXDl527PrZiNOLJbfJkkK4TRZF58M+aAU8q2vCI7OMR92x+lTUSIQZNB+
FsR5M+6OCT/tDy+NW7oKuYmBgOHIIogD16RCOjbbGecIj1qf27yGYbAPiTidvcaz
apjMZf4yhKZVbiaAjLBLQoDg+1mqQy2uqgOuObl64QWL9eCEi7bC4Vtaq+acQ/z6
R3W1l6Rli6hTlAGbdSSBr0kykeFJjnjVAPSQta0o2VQQ8OYWmFF0Wj/ZmvVhRAMM
aIDgwvBNn5nmIrHzpGWJ7ZxvqKHJFm2+3YYOSQ8e4F6WrW6WPuMR39ud/3zPDU0v
WNxaan7+KNSU8m4YUu5/7yB11+2c2CheQhhdJwsMM2mDgTAK3M0PQwAB8aD9QLjD
m5sm5cFKpQu8RZCFgb3rU/FfAFuBzZHPzsbF/f03V3Sczl6a0IKbcqTvhcGHAW3+
ySquh37CAlj68p9TeFeNNNF2OXBJleb5TZ2uy7BW+H3w0RsEwQYb4C21+IAMegE7
WMDNnivbCLsPpPGwohnOSPkZLwSjxma7antQWnxym5fKfgltMzNHBO5mL8r0vG8l
rgn/PISAvMmv7Unlvulx2eg9re3lVojo6Z1+NVbBelwwXFwGQESAnslxv7PZYRHC
nxZRAmZ4N4bFep/rPpOc4CZQcucC1nvZ14s6nJKd9Llcqrn0By/nHNyRNEtRkJHD
XjMfqN5G2LQfG9NMXm80X4DoKMHkAaw4VkXAOOR6XjaAzrDPsZscg6rRZD+a45r7
42ZeVlZeRcdT31K+rwvYUWCmp3zO5jSCSog05INWuVBlKxc3ha/GPF/dHEspCkbn
fzsFg2CuLpmHGOm1s2l4LaL+dM+29QnxXYxPFwao/vkmBRef/hFCNnSzGZrkYPye
GXbgCotQrPFT1TOqiSDCUrIYPqaQTptK83ny5RtLybG4MyVfd4AmaaW59sOgZQDH
bhAydT9RXHXYNqqSZR54NQtu1unkNvwHiXDmhRkTv2Pl16yJnpGmHqkd0ZT2VZy3
o8lCUDas1O6iGrC3nEXekMoqlIHnE4Kvf9VlqztM18B8EV8RhUk2SulqAC4YQ3Om
LpXqLjA/heYAY0thdE6X22EhhBV7Oj3KbF+ep9A2U19iiNTOb7jp/f6UP7GuS1tl
rj4oz0sNoTYcBuXTMzhyoY46Ai2I0iYZ5dni+0QhoKC2YDv7D7Nz2Q09j3mI5TtC
CDpxI/zXmK1s8lLeIuqS6xagrsP10KCrKTmtggpAX8XYIA4mZSnlGsd0obUTBnAz
vsG5mWzJANbgx+az3/ZUF1V4CjTVqPg7s/MqK1gcYkSHS4hlvyrxPkvqXfgSjP//
nICAOOa5XnOaR+Vj+KMQae/U4yedxTlEYw+N0oC7qxdPMOpCYsUIe1ZHAoV936JU
lHqM+6d8Q5aQg+kOI9mV+VK+RTEjg2+hYbQxiFg+S5CcFztd42ysZY0Tp4+WlwYf
7cWOX/4GCHhuKAJnj1BRe2Zf3dRUYJiRqUhr5gZN3PUpZ5bfMtHj8z0KAhk6g6dJ
6OgsZvMAMPh7iURv1sCiBZOCaBscp8b6k/DCZEgLDJW1r7SmpnxF0zTwXpxnFo3J
rvn7ONq2N6OAuh0l7HtylSYDwBw1F//MjE7H0emFxF7eZ4O9ifNdJd/PTtuAEe7c
692gzr8erkPQ3sMxXV34NvSvk8z7ynLbe3jDk30/Vd9UhW/xe1FHDYvpvUfTq+4q
hT0GXf6VYwE82uHpYq8xksBJPRh1rp6c4vdFXW1Zw+qMSRU/GOr96xccU2Hoh8nY
wTqMkEhGvrnhcFfJss8kQE2IqYxGoXDnTWCNkTOMkIh1DVcyn5S7GttwBNhlEdbc
jwI5xhZ7QXoMYV8ihH0jYQdmoujEkl47BH978Ow6xcJW/Is6QHpf9b0WfXub/1Ok
GpAjZbpLUbwXqWeYptQS8waKbRRq7rlVOuLmHtYEU8o8t1LFcej4UZOhfzctTPVh
Xefh+B15Egw67G3WrQJhwnuGKgb7TXwmsGqlgRItLCC2I79lHrAvbuSWaPBXRo1I
6phyGh0FsvVHqUrkM8ua4vnUK4IlMltjC52db5HGMYrOqATLozetHOur9qlDEknW
KOsa8c7jp/ygg5zajbeWiyZmI/qgw4XHDw/8mT2ldwqKO+glthPYJ77Fdmimlw/j
Jj6yMHKaydRz4mHdDaz8g/eDlytOzmZ04vTX1fwCSdor001z7t04bJFg3wTIw1ZT
vcj2KjjVuIXqYCTKaAIDvO4S7aAhKZ/2iItWw81BR4VVH6BxQyTsicXrSESqRugN
P+esKzZkPXf9FOzrNh9aDp66OPz+RS0owQ5mtMqcbmYOfeKqR2wY97wCcWEfQLA9
JsStu/tkdp+uUMCY4BG6JgXHs01XDGMy+tb1Kfvz+jMBWL6bECmZ3kMJJoH7p2O8
D17Wy1rVrwDFgwQ+XaQZKNTVwxyEdg0+YMkaTv+JOf0yWFvXtxu8URAcP1UVi2i3
4isQnAluYMZgqal1rKSpmitNBshv/vK3PH9mXdBLM+Bp5dZY10KMVy92vT5PEG9N
utEj1/CKxicv0o1t3a1CwoFlOsDIjr/vq1SGrCGMHlLkBIxwMqxUPL8M99sEIBeF
+WOQpJyPmt2h8hYWl7PHl/yQZ6UFq+Zy9sM6FgyOYb83GLEsngQVGhBVge4g5aUK
CSmm4ZKghLDPhNVg/5E+76flg7RXVSi6LQPR9HgFUa7H74jGAnohBZoINIGVwSFc
weuymaKNsEfps3jtXKyGU5gscpdtsc+Fqv3RKUaLAamaMB2cSWg7I6yEUynp1DRN
l7o8sGZRy0+oZZ127EBG5oumT5fnOJErAea7LVk6yeT0DGphZaJGQUIdXSS85EnN
nyDW0G+QkN6pRi8VoA+XDoKiNo0SDQPuqGhUTtj019gofHbMJd3AokxI015XAxON
JMJimCbEtuxaYj0kxlSal98wyB3yVw3VSlhH3cHpCU0BYqILvRXCr7Z2B5hwcPXL
DP6G1VUFvVYX4/tP3UAcsYO/ZI3CGWnmJSZC9moaobpXXfPHLs84L5YQGJdaebDw
Njnw/bDTw9nM2rc4eoI3u17cS4oclucies6L/OkU81k14/K7HrEwv8zZ9iEjMMUw
vbEQSkZFWqiZlyJoLT9AJCznR+JWnpU5jIAJG1V9udDBY6+5lsMtXqaAtitckOgY
vz20PklwIzZTv68YyN/pcI+MIxiWRpdLMzL/xHQ/RbsKnotMF8MmZrAyiylLAvkG
y9H4hWJB4JKk/7OWPxDyn6Fxw9yIJKBn0zPzTTTNUZR8wgdyfWtjK32rp71hWqTR
vQKFgzJ/J4+de/XcLLnzVU1R4h2HjS7HuG+qC7L+OcQn7Q4Omg8SSHysj8pH+9FM
1Hdpg3dz2/RhHvXckurhvm5YI8cznYsuOtFrkvltca3OqBZ+Mza/z4t6ZsWFvWKh
VZYcGXzKdskXzLSrr7ymGSKL9pqJ6wJzR88AhDkumgXkz56wCc+AtLgaioTsWYIn
U+gXHAVWUoTHpW523IoH9HV2dVJ+rMhOKwlmEkFCarwLbOIJ2sHl99I/XtCJNAJU
UWPStFrByKp2a5rW3JSYkTUxQeyE4/1qm+guhlTb6WYY8WjS3L9/0hPQU34JpmeV
qYJ6siKohm8sr+pdWkAxmLl6R+3QZtHIhg3g6Y59HR5kydHJdqyQnPyy98yy7f4P
WgZhqg0/WP8P6RipJSQm1oX1ym3dWrcxdksMVaGKq5eAWWyhXMjklXHTj/vluPEx
6sQTfCM+6seQQeHheebH5PWQbJVgMB/zk/Ox8+anE0zkw7SU8Pd9aI1wiu0j8VV2
xtPjZIGvwRVLVEXa/bJrbV1jo2DcXtYe25LG1XnKK1dk03DaAYqEpE7io0F8s+f8
1CYKPhBFJaeELDY4hke9dC0yqAE67sUu/5kCR5T4zQHw2E7eunIUGkk013A8T+Py
l56Qjra48ep3ejBNdoYRX+e2IwvI4o8RspNHX4YtoGOLi7PKDKnCx1v9OArsnRqt
Yrmp8K82HVa5aSF7TKUEZUvJ5lJtuzbuiG8/XvJGv/9ZUnhSdI+5wNf44uz+0D5+
/1CEkX0VngKYbQlBhXEU0YAeEIiv+CKGhdfWqVBEb7253ImwSbMgRYIfNaZPImVM
EuuR9kG3LCJyvNAYmk/ICI/UJwK8H2DtIFCs8CNL3YN5cfjCLNudTP9wcSA9g2AQ
jgwPTw9FPuKzeTyNrtuJPStIc43EAnWIOyECgQHSYu7ogvCHKGRD6Z/rMnTjfIS+
Y0X0mRt4eZB5MvljQNAqyhQzvtnLCsxAm9FYrx80kZfSP/sQcXyyJtTbWkIeKoWd
uvZdhpbv/ogpbcAkQn7ImchepF6ZejL02dTjtV6jyVXPnDJsoRoYCiwUGXvbJDfQ
hlqw1p3pspPt+IJQ2yudJg/XWojwSweYJTcyv5zzQCcdueGwPccvFk3BkfJj8biC
rubPYReK6Bsjky/XTzzSy0ge0SWBPQVVP5EfwLYcmPZ0kDO6GnHhV08aXqw2iU+T
yOlA+ARjJnVYdhG+h2q2rsvgFmgbVEa9KaoF54g8z4Voy7GxNPGmUdlD7FASVlt8
IYSd+s9BJ6xWVgWV/32KrRseibORr0gEEkdeY+zGfv5ZSD+uCqdC94Kc9GkIEdPQ
6Q6lBpBZv8nupcyB3YxmfVA53GEYbmQmD5Iof0AvEf7wnNYgVrny9bH5iPTSniJo
53h6dRBrMwXMljhOnUOpbub+IroCycnTvEYDgz6CuyBifrxK41GPe32PE8JQXgsO
3PJb2GpeuetMmXdQF2OIBlYYdWaASkIuGlKogr/eZ8D4RGimPb0suhjA1jjajDg9
xXm5nBJNleRPNZqwEVM+7tUlAkWbCDtFg8MTXm/bo1QdBBgeZaSv+TQIFx343Y/x
bmUPSIldnwG2+9ldi+MjOARiDnhTnXVJTTwcj1vjZvSoq9N4QzglYeqdRtJVg4Fb
bYol4rWzFMe3PX5k1YHgl02gLn7SXXmcJPesGvRv8t84MrPImtCYFQADDK7qEM/9
lQAySYn28KrkOX7+3Fu4nnY6oD+8TwcQb4moLw19pOZKy9ssNdZ3O1UV6MkeKrkz
zYSDMr3jGhhM1BEA56Dl+R3UhieTnBoKDmQSisnkyIvARRZ5zFVvifmz4Nx/MSVw
vG+ImaAN7wQHa3BPVEvQ3koSUT5DW3JzY6LfPdCIZcnkSjS8PCPeJala2Dr8Utlw
pT0wyViN0njbET1vnddVoi0Z0qoLCku/tG/aIYVio8N5ZFMUq3jLwgBqmSY4izX1
+vuYiSC6KNQ4U7u2k0a7yGAPZbem0ND3otwHoVvXnheJHDdEPICc1piFQI+UMrUt
5koUMvNd0Ai9lrA7JOwh47maI6aiySkHqZXWinW1/7DIJ6tFSufDIPWyWp9mwV8n
Th8e4odAaxU+18lc+9iptVBSI5ZdW3nvRVgdIXRynSsuGi2MCoDfhv6jfrt8OKyF
oCVZqC2aUCFwJPf2ft4b0IJJKZ+YMPchx6aWEEY7V0lRueYinNYWsQkdJQpdJlk1
zgDNoirUXZNBCrO+8rBZAfavVT9NsUCQVYrKbIGVqn3HhfVvtk/ZL3A5vSnXkwZn
3DGZOgH1MQv+giesg6bJg7Uyh/tITG0NunLHZvVw4G/IQVII930ajmKhZ2v+v0D9
7u3R+iwzqhRhFoi/MS8HleyK+aE2L1PIgD7LucqfqbBetdg3jk3F+0Hxuf3e2UkK
+AZNeC3v6Qf7QDyQquPUaSsCNS4Mk9+CaWtdPw3XZFflnToYvjo2ppWq8ViqVW45
zp4ZDbTRZELY5Hzs1LwUAMgTBuupnfd3VROaB6/Jw0g+BI9Dmh6mEkxFBaTY+pKW
lSC028aZaeEHX2jBDkZ0ePoLZTQNEllO6zvKmL3kCHKxkUMV+hZWXmUVyIxMjTuT
wLyIekjCy5pdW3t1XJlAeXhOQCRYwcpX2LhjFD4bT2gh+hpMYzpUrM1o6A2MIW0D
3usHOdfbVou8ubkZniqCbIxDWLoaECDJobyl+bsrVyxLJR8atd2wzzakNbmR02xl
b3oymx01trsXVrMhR2poI4W/1Jx0rfEe1a5Ov4h75AzIoRIqBr0SKMGIpYkaTyUV
Q6c8tLl0cM3djt20K7ZuhypcWmnje3ezexm/xP1fzr4mHcnyxAlsrd0ceq+kUclr
qr5oN891ZwQDJN22EMSK2yeO0hV+F+ZpeKTq5IUduqqXjqD6dtZ3ePg/gZoVnxT4
NWP8RzCWz1WXY4+ZbP72oBhLH+TeNsKWzeE9goU7cd3BoOfJPbMk1ssMOdjrju5m
Kpskw9y9a54U6kzETfwdcWn3mrQH0N3kjfFt75e9UWqffcB3vgkienK60WjyllLp
2M3WB77shiKVNw0n9uE0cp3aXeUZ//S5huqNzp4gVScK3sOJxX3eWbfvSOOu9v25
4L75f/j35afA6whDUHT3RXz5H2Q2q/ahiD4JiraeVtXp96WnJQOjYVrIhrwW7LpM
ULEZWFptAbGptB9+/dF2FYWitDEftFMiT4+d0BmRSnyVyXqemVXjb3LFAIqjGTzx
mbvLlsngsic7SYZKPsik+IRuwwaPGSAlv2aEitSoA8SK5UmEM8J8yHunUXh+LEn6
LYtsvVCS1f5GWXg4GrCA/OSqeCuBve36aH9e9w1FozuXsWCOewyzWTppD+iOjgbA
j3chKUFtqar8Hnuy48G5Al7XnyHIf2dSY2f0jdKkiUirgwEd1is3yE1JQ7BlF6KH
oftQg0EWGkA5gJrWjPD13EvgJSYJ/jprQ8KGAAwzy+0wMc/U2jTt14U/w6TyG8M0
SA7MhbKwXdB8qjadoUqAuoPjjjnT/LM4FJzmI/zaUOOyqSFladioZl80jXpvZ79k
0/dP3oOnUJ5pQt3Sfopoh323kKj7rEBcIaOqtwG5g//gbYOpzEA/sVcVc4+WZysc
83D2IgfdEh4ytMx6ixLcwB0Pz0QIW+whNPXaUfzdvc8Jv5/mW/zCLshezAWZQTa6
3N5PL5Y+sWbZIVnG+Dhv5a40E3XWure7JdFoRRl73kfH6Y5FWbofJ8/Wrq8KyAz8
1jeHaR0IiQtft1YH6xsWAoMRyNKlCw3SP+7xQiEN10iTlppBcLhe5cd4VF1Pzuuq
1nGcle01x+KMqFLCw4xPggh3fGQ1TvT4jkZwTyHYy37Tr4H/myjTluj/KOYjxvL/
15/MtzH1e3iUBR+kkzaeBDLMTFOUD049VxYtewcMTF2aJK2gQiMqFllyaJFtRLM7
N9IJe1S4ZfNDlfI0ns1A6PUQUPilDYp4SzwWEztgDe9WQBXPYXC+fyDgQN9zvyY5
8tZjfkqzOoinBav/dFKS/wwzBF9zZSme1cTJso0j9dQAorjwMfOWZ7F8vSYN4QxC
dXrERkDTTYp/fpf/JDjtiTlY9rwiSWa6ZGXBa3rv7Kyy/RKBM4pyXd8xe1vFh45c
JH/iyb1xuwD+KsXec3siYZIPGXbJRMIplEZ019sRAZivrRNQx8k4DwHtvfJfMKc2
I3Net6BkSl84MGJ6k8PjZduCURlG2/ySjtkwgODnQ/+HzqhUOzrXLNoFfuSDOrNR
UEQMkz3z3mKBVfaywjixUZQFKcRgmkex34jtBi4B/J9JwLqaQOgu10Qntmbe//r2
RwJcjQri82qhKED5teui8U5466qajgVdaIfzxVwy4J/+TXl9L/X+0dn50+ShPBnA
fCYt8nx2YGndtRxnNFFZD8ynyhGi56JORi4PfEi79nQ65HILS986FAbjgj2zUxdb
9avbhdO6Omq3JL5XhTBUuLuMeIYTrI1lbC5wEdscoM65qq164XtyJljy1thkjzms
ChqmPXUGItHKGV9fBDDSmfofDRlKhDhA26UAMF/O0BmvI53X359kgzHwZO7uHzMw
GKE0VWS5F8k7vXp962CfLmvesJNZxP7IwxO/waJ5ZGzUA/Ev8r9GhKbw/H83Pqen
f8YycOdfhZXP3j7eQLjxvguU6Zp8FdqHxj6SLVeowIU9sFrDNG98XmFzRpOwZsi1
P8AZhwkrTRtBD/dEvMJS6jwGKSYJRkBNRIHpZftwUFB4mdTJ9pZqgPp3Jt4SjtDs
3m+iBkMb1dS9oHpjCUPjgUxqLwAIzwgtPj6GSsUZ0zNAoO64nTTQSUCvx89lYc4J
Qia06r6qewX0cZzibhT2D/xsOlxQhE5qcGRdBYCW+mQpLsYY4FYVe618hx3D5v7v
p2pEKVpKQ0BPV35+vEHubithfabDkxDaj/xT36IX7WmrC/pHSiV3kqifv3MycN9i
Gx21tez8w+nyrO3YSKSh19Kh+qXZa/0/RY2lVAC0KHK6iCRI2nFGNLzzFkzxaG49
ailm0UdhW/izDPgoWlaw3q+uA59UBDmCT7WkKjrQDLFK4LeKfrchOtxpwXVyCk/v
BELUDxT0Q433aU7E9lI7+KmUcGsVe5zXjcCU26E1gOhpzMLE1Od57aOEWBP1rCNS
0U0ZJKYM0vyolc/1B+FU4kgrxpz40xdh9CTcRHzw9Hr70JIOEPfTlPM0UPVyZ+er
ldsK5SoiGBd7d8oA9jr8DQUl5k6OL/27McFv2NWazIXgL6cVyY2qbOjagfuHHjMY
d7KNhjGUsxVyU/ElKD98a7M+4NXj/VgoIA4Hmv5tKcYH+yC1tg7ScWgmMewCNx03
2xcYgvaC38lFrMMmQm14hh5b/xCusAdHunfDsNL9bfcoJH2q6KeBUh0g9wnQ2SHk
qRM7hgR8hW/zHb+bjXTJv5PjFFGoeIV3aUrIP69cf6D/sxwSy04tuVIOkh21iFne
0Pkmc1YfsSu3TRtASwg7SoBGGMO5aXlaWEva+2ArY1S7wx6aehWXN8C8pSFw4CQE
6CPIBoLxprVE6sfWe6e4vG2e4GXuvSsDJmtx6fu5Ozkd6PO0xc0jJLc50NcxrF7J
kZMOE+/JVNSkza6fxHGllzp97V50+6OPeHkELP1n/lxxca8zJcdj5jhMgkndPrn/
h037PcLe22N5O/xs6RpeeFpgqOXm2iUaa9CAELR6sEP2JiYorLWox08zPqaiDCAb
neZllEJ3elkfob9badUwvxH90DBn7BMaqklNFAV8vLZyesr8lpFaOUZCPeCGcEVI
3Elzw20AgpJNT570WNjutxrCqTgqJx0BpvQRL/S6hTGFrd+RrEhh0/vym+uZPHpG
TvZdqVKN28scvoCauVaNcK7I8ESuQ41SUoVElhKg2yVrEXlmn3+tEYcU4zV2iGKh
sFy3nYgWvpv11PslPfkGE/2u1HfTMSB3Ln6wMeG9Rvgjni5j0hCbhvct8QcH8/1j
1o/QPMmjMGOQiXNWPXbAtIBBqeSPNxLc6C+cnB3ZmoNguKxatAsUiaztxaEr5gTn
2o3PICz2A4+H36FTs6Oknx/heyMTRosLcRCW0rg33pSGmmVNgYWk1UOBIXAKhHwo
y7wpAondKm4PCUXTdaDfPI5t0ecCP+Qkm8cyoTnhQ/+RPZQ8F7grCwsd3G4Xkse1
ftUzwTyyr0jI4it7xFXu5hjbaHp/8d/hjtFUJCrNoWmpdwOFGyB1hCUo0IXiKa7c
1n3ka/iUZIIXoel0yIMXx9+wxuvUw6DJdHYXqKCOtJx0HLkKWw5sfTcdDnRV4sJ8
VGx2lfs7hghQKr46ZFYKn/N39/xsJrdxIAakSN2CoNyqMN7oEXeM66WsAH78bohY
rX6XvGdaKfqUEKyBz5Ukhsp/9Vbsw7j2zeJ+rAaztD8yHql72Qz1Cmey8SY6gFSA
WyCdQCdwPFAilc0JAwVJP6ZT5SDzO5S9wzlfFOe7BaDGGCMCiKb4BQrOHycRITEU
NbMT1g67G9CpOvV4fV/gzOO9ofptPcalEB4mmpMhyhwryqxrRsmjd8tNQKX7hQue
Xaca1MIceCbXA9jE1P9/G9g3VKZwt9/1h7Z208wBlg8BJyzRuQ7tncjKbjIerfRs
6G/nuHOJdtkqrYJhws4bddO4GjGxfqENfuFLPg/stRvbK+JXlyQK1s0DgOOLr3l9
lZx7Tto1sDo3vBfCPT4QmXZoAfA24xUR1IsXRfYTXlNu6NbVLvCrpuP5QjU17Rf+
rI0mk/7YDXw7QDDaPnpvuXNS4GY7mePnhknN8MyHPCOPKnAseDaJJLpdCxrbPIMm
aNaRMdt1XexA56/qIA0m6HafXBVCbaxlC95NDnJZUFzxBQsmr2ITDGKzq+7lu35F
FhdUEMctvtN4sdk/vbKKjTIhHZOnhCgfgbQ7Apngz1WntpMRr0qpfARdKU3Sxidu
4YFGlSU1apesTlfPxAqVMpBJAVXeVt24qHKjOtdWvj6o93rHRUddvhzjSegg6wmQ
UFzm59GgpYu6QADBSCFeY4BEtxSFtyc5sRc98YBYZ9V08aEpMxxfsc45wh/XzaR4
LhidBJGtEAKcSmf+PBKrDLKiE7vEWFGq6LY4D2580mib/FS4Hkn7haD4qxR46GMC
rDCasXHTnVPG0UY6sg4uA+WTgzxIszxOtZwDdrrxgIipQBx9U0pCGHnHWI3GRWSd
cF30zJVVOy1R3CZp3AxWNS6pbFPKxDX1PpoI6gQwVkr96p77Zct300BAaS+V6CGX
uT36L9SePqCSJeXa9BPlvpsxvnCGR0hWHOfFL7CkuobxY9FIaMaWY2MXkMMwxqCA
rhS+8PbCKpTGciJbD6Lv17GFIwGSf2aSRJ6d3HqWRuSfXpmMYXDrqSmihnZJhohP
3kmJnXvBVvsbuyvP6WDBCJVjI0eWOcsGN6EyY1aIgjA1vGLKcKp769vGtiiKcVGi
1qkszdkCkf6//GoXPaQNnFgQqvqzZ1VSttAEWeGw4XiLc3zodAn9kX3vkbYkKmfl
txGDhg7Wz52Y/+hZqqen3TvybjY6FU/EbJ31H93Ik1bU7zolfDQFYiK/v2svE9kN
sRdg16vRjXiV5ygOIZpSz7ix2mU7Gi45hQQ/LELzR1xh5LsVpVc6LdHI3+rAaUzX
fRAtUjHdCZSrNQTGGoJgcvx0VqqBJfjpiw+gSTvqWyAYAy2mlf+dkraEdTAyAIwk
7N1cKGX6Aio5EjITPI4swaVXwMEI7CRQ1xHt/z4xF9PL1xXLzQwQx22Yl/EW3hKx
OPd+0nU1gfyWddBeui26XrtDWucwTy4/VFWrtLXy+tT2zM/9N3RIqN1utTnVo8cy
17nUk+52UNrXojbf+JhEzQDcJ/bHW8h5YHdeFM1CN8lnwl22yTXiCAgjFbGYKS3Y
+FAm3Sr+YwIk2FwJkleLq+NrV9CYTc82NfIswZ3Co1NrAkSa6N9f0wF+Tq80EWku
Hvltvu1MW4/BvdXfAPMRweGDE8OBpZHJt//Z/gEcctUMengJ9oM8ft1zwV0tLdx3
sixOUMk4/P+vkUMdhoJk1tO7Ujx1qKiAgEG9XaO9XqVbeu0CjvBxnLaEkJgnc2Fk
rJi0xLzVexHQg1u0ZvhHonNTmeSPW6ZebYeIkg+irBHCJgHUWrYWQM7c62Lbk5s7
pJJlMJ5mTHKRR3Hcoh3LdOC4ajoRytN/uNYRZFNWTln+w8g3tHWCx/IRlQgpPnnZ
39zv/ReC0uTGm36Fs4NFclueZ61ptrlX9QFiGj0WFwy2TV1QlihYzItytqV0GvJR
QD56BY4r9JRyZN4KyyncsUzmg3hqLzGghl3KLZ/HY7/OgDBCgQuqpyp9ZmASWAx7
SL2T0rc40o9fqrLSbqd03YkcYZjXHSmR4yGGpTg0OV5W7X0judGK2Osjt/5o/Fxf
WoTqegUZS12vPNb1ESup1Sm3xce9hnd1ldHfGTrtCI+pTnfJTa3ObJlUCdb3T8Ja
RPxBiIL+TqcsWNLygOgVMp/P2Fp5/iKxm5WB5MMGmPG2SBJUYJEajJlFwJl9NXBu
eG2iaF5CA7ErrwR/VmkbWIAIhgVeyJGm+vcqE/FeZAucmdNLyRhIV+3Q9XGwOItp
qmFP4pEs/DQvhi5x5iYNf/hq531Afla5Ysu02kjy02iIiGBy+UUqnSvTJ9IDB1Fn
/XkopxVGVP4NJ4H0WIBdUK4zaKUtJ1CW0B45TnSJC25ZFYV2UTgsN/Qvc/2QBYkL
cw2C4Dby8PgTPsym69//Uj2gpsJLgnoaCS4LiXG/ZDuTlxnXPchcKQnK1cCqF32W
GCpcSp8LR2U/M1bE+5YrYf3URTGLlhkdn+b8XDD3TO7onIhq2TEodXyIpDJMaTH1
ODnFm3vOZMs/4GetAJ8xYfxn7MN0kVwkjcuvJAbx7Xeq19vp2gsg7sCPeZW+3nLX
CIMuj/H23FB05jUf8W/SMK711/Uov5Jb47gJBL+HboIiQFNm7hCBLZTsusXyAPtB
i7jHFB3fgfa8NEX4uTjlxKszq8ilxqUemacTUnU0FxwxgMdZAWnELjx0z9afK4vV
q1rZkpmrzfTQR7wmlV6BPnfsC7ZjBIyLbc60xSt2jKIcfELRmuhQhYaMo2Ho66HZ
0zg1W8Kn2e4Hd6P0Rs4TfKzm/c4V9NVu6dbMIjrAwyGlLOLZaKCa33NDBFDNYMZ1
+d2k2C6tVtHyKpdUmDAtgrGR4i4EiUQHs4FvgJR+b7gzKrZwGvi3fcVpm/WObqRf
ok8m761zZ40P1K7svMLjT6XFo9rUxOgK9SOPR9p7DXq933cluLooZ6t5ClaXXYRK
6sS7G5LM1kJ413mHUmwrTW9uFbUQiQIErMiCEbcYC3mfcW+FRGiCpqmH0w5QbzCg
5uXmeslLRaydSn+i3BYAuq3RqvXetGxAfHOJOxH7EqHJA+ZeENpbegCW4kVbGtjt
ehdqdcWBMCLbqtiNYmUjGpzNdwzsOUpXYXMUTdTRyYMLi2l5ymDNuZH5Qp5q2sm9
URdsLZ8UQAnwazxUT5+71DmgQAaWQqLLvtBrmhhc8swdKKHhPi6gPQBxtUJqdwwb
r4g6ecrUmUZhR1fbiW7NKtygoDIZTDvjE0mHVAHsbpasYD8goh3lpCetmggQDpXF
AiX1hEl5a0+c6CKYj/3pjTDrccjFOoU+UNfg6EdQAfRMhzeeQbwPyW6pinnGkfjp
IfWW2EXgE/eeIpqV72oQ8iOtQC2cVXYfc7idxmMn0Np0XkBXxcqHv5PrdaYEnJvw
aG5EqLxOlJIzyxqxBgoAQ6rylIRwgGMZKX4KGvH8OJeGXgD4Rc1eg27atjPURigM
YyPYkjjmGb5eRJEVVcbcfbml04Wrsg+girBC64ssDaTDu2kjiaPPv1X7alRsqRo0
O7cih2+eM7bjc3zpX4hIgHmpcTcDgyQSQRM6vduzf0soG0dCwr0HTp8X9FDX8nof
KKaHATRaOwKpTRI+EWdjh/o+gVPgdLRa77vDnoFRu8K0nBZvTB4AIsd7+zd5OHHa
5wilnEhvT90ZvGWUt+PNzsEtKrob09WDuUFyEFx3V7Tq1y0bjf20L/yGwZf6iQ1I
6XDeyXFSbtgsT0QNJ9N5wdrfp0Eu3X7f0AC3XujcMBxbv/zNNwW+KoYIPlN8K9Jd
d64MlNSZpyq8qV78R8DY2wTq1YzPmTTSfODZ2adwMFLuleqXw8+tHe10RXNB3GsA
o+DmeM/T2dYySpaIATkCLNQ7SuzP+cKmMKjXDNGkiwua3LZhTt782YTVXXuuasFs
Su0tztquB3sEc2qkte0wmzb7BpCkZTAOHG6TUYMRkCIWPiudUI0onmUB58HMl5wG
WwLSVtuX1EHIN0tU/KqrxCfXfIt9FuOnROYDUXHmSFZ9zsFjnKUSecZTa7+EXY84
DI51IoJs+OJmwk9Uw3w89X3s841gKpOq8u9hOtMdQ+f5sq01OErj6Bch2y4G802p
6C0grmr6otRwdz9pV3mgIAV7Yr+swt5v3LuH0jHcL+x0nW3aKdhHPPj3H84UCEEn
LJ3oH0YZU1KnHz2oQDD3W0FeU+W5crHRV9Jbk5H2IzWS0PZGWzjtmI8mIGdVVage
LT34VKJQ1esmlnMHNsgW2+eYjurmfef4FHj3cqNo4TTCdc9jcCF8QpIWdW9ZZk4o
6aNkDLcx2h/EpYd1oY34py5LkgbGunfGUPH9V9g1uKBstVEaz1bqZTHt4w3BFyY8
8BaQCXOqC3WMeDt19VrS5zqHae9hJ1qb5GRSxCF4n9StkFkw6IEYFwuY1uLYF7HN
LzLXJoXSZyOgOjzD93QO3tHf9pOdVSGM+czjybLrS+EEYWSv6ybwn5zWlNX8njiq
k8BXzHMSP4V3osVIqTMGYl3aEvX7N4mrqHaTEj4k4ZYciYJrWaFsv3M/IDgAJ5T6
gkfVwEVvCLXG0otl61/+yVAJZRf405kdOw8BlZJRGYuNMhgaTCeaG1wCqzuNa/e2
xiRLwJlKVCJ+IIRcKgy39nu36Syk2EsSMt6Fv6/enHApzUsnRpTI6PC5gpIcOy6Q
2+Powcf8E/6AIoLLPQhrXyeAo0pC5tkWSOjQQATChc5Q6yYttFYiOC2SbpiZlUEe
+PgfSLfx9Wb0I81B41yEm5x1SffiWD7AUJFUITbCHZS+B3b57B7MSJk83+WELzi3
1W+qDOPSf9ekpUc7EpwDyI7NAcCOUnrrJ5s6ZGf5cuX4Mxz76WKtM2tmj7dBdaFx
mhFKSZIROo1sJZrXS0mWOWeLnPrEu+ea5fsvs8k6Ff0EBEdQ4aaWLmOd0zV8XVoU
kcrJOkfT5FKHVZTWOz6G7H+cj3amCvRuVvq87tLbeA8py39wp3jTppyGs3BTnIIT
AKY9hW0J/HykQPT889suz1n2Jh4hTqY1uwBOMjC6aOHDVTbd+fTdVcz5OPii5XRn
k4ll7mOBONiA0z4X35rL2z7oYEJjpzp/FBPcfV/R8keZ0n6HABmmVpQx/7lDKVMm
d6HVxji/2wx1Iv3Zo3bkKsYwaOr7yFz2fewcqednmW4FnVjzCj5iYHmTCmInkwEu
iZt0CxcFdJKxGHIVRVEtoBtViW33L6kDdy2xyaCteb8TJrNdB3MregrVX1CAA9NE
otHpDKAoBLn9fJfQsZljxsxLq0ERBNo9YwYHh5rcTbJ7x182rEnBWLr83WvkKwW3
A8pJpheholY1HF0qMmOoJ3S+qh/spKm2HtvRIjlcUxxO1ueBDzc3SkDFRgVODdqp
fijVw/kz4oGa54T9nUKj3irwK1zAD8B7dSXW9/WzDVImaIt365g2gEgQLbUAfyEK
e2GcF/l6ARjX0uTaJQPXfcASOqvuPwlAk1JuAahPfY45VAbj3S/pm9+n5fCpuKoa
lqOb1zdXYJCKV3AcXiuloo+zCwAjXLjWpiPIVhcvLVm2eJufrqeKexRo0vRD5dHp
Mp8xKJqCWsQeUJEbAe4JOQ38J6TWzntUA2syPzSrLDN4N9lpVMEtjHgqZPUMvBcx
Kfn9puJqbpXGAbWTon+nBOLVjUxPZg6cb9xdtPYBlJk9UPBU/QIvDACJb7PkYFtp
ulmUpB9VNln0WEt7slbRZY5j7j3zNhojBTycmRxoOHNCJKAaMbp04h+1yfg0ffX8
A1Y0bejG7h+i041njoxSZ7bV6BzhTqjLx8wfPke4hg+7VFqaU7va1jZzC4EPzAqj
+8LBMfpcaLnGKq1btSH16aE+armX0ebRbSDibJoEYzLA2lCBDticgxHCehPdcFzc
IGHxchNRjeN9ZZSXLiBsh3z7gSfgp5NOf+RQihLjQkccmYm8F8k2wxZ9rMqdgq+R
nh+ILn/dP1LzNTHwr+BN6q4WJeZoLucbK4LOFj+TWSZtEQFPDFFmcfpMhiwRL5Zw
/iqJOeP5VTEP0jOb9Eza5oiUQSie+NO/+02f+3D8LmFWTVl+ou3Gl085kSfCvfcn
dYK6fQuANr1vhRvz37Yqdl4T6lcj0z9jdKMa4OwsAIzsJotPyE9q+sDnr85Z7Ou4
fp1Yh/Coa8ZPG5/3+DFQyPkMTHPOM/bA0gOlxub3f/uKg1eKsrbfVsln3wQKW1PV
BgBa0djAx22pQOBcoRhQGyK/GUHu5E9ICu21PCAstozBREF3NR121+qYIWoPAS/S
sWKDEzn6YrK2WT6KijChsYVXSzZy+c1JcHwdmUzDopL893zXrWOvPejxyxcuO0I+
dv4Mi/gsDLpSC49K6EiaMuSMUnhtuIpV9EtQaW6Joed0SCJ3M8OBGjSqIEwyHth6
BFEjCbbsmpIgITz8c7C6V/W9USVhhjrHJB2FszJE0qOLnhDEzQKQObHu8wDI9QQW
4vmNH4kGoaU59+J+GuWr6SIcSIc/Ju9AwrCEoqzQ4Q0VVL7wrVyB/su9tme5bKFj
JjyEzPprScAWHll4MqAVBvCwGEAufFTvrZ/dCZmtMJojYYWhPvaodRZGHBreVEpf
kDKO9RZ2z95xBJ2xuiaCsy07Sk85r0fOvFGMPMxI843hEnDsvYnvVo0UKVjSEnus
M/8Bb3LLqPyIvGDYxiF+SGqAm0CLnnlvEj2nIUwZYF53GAzBpG+r4Vy/1+I/tQXE
CHjf7DjbOl6WVAuX51jPAKa2LWRvCQrn6jCaBYhne7vIyQ5nfInDY/QpaXWyO7iV
1HZqYP4/VmWwtNRlZsGBtUT2CCn6hcFKywjKm/WoN2N7T7WPRoSbtVOOHoWZMguG
j9yf3KetdyTB7nv40PBGCkc0TtOKT9rIcI0p47sBKQowIt0M9pUrZOUok6O6Qqfx
YwVQS70KtyInPLtc2H2Vtts9gTMI3JPO9MsGh8fHAsl6hNhPKq35QzNSqTHF3lnL
HNM1ngl6feXVwlH7i+DIUU0Eu/tcb1JC50luCSsl7r+ajemEgqRN8wfNcQKLvNlU
GPaIZIb4e2Cm+ePhpHCNK1EK0Gu7uTSLNqmf2LnluhOn9/dBLgSfegpxQiykF060
eEO7n5gBnwSYeyfrr7H0vZN87SMWv3gTUJ6IwT7prgkILAIPocu9lHoK02trs4gs
GLN1hhB6XeTjKF6fo8BDinVCRdA6wbThMeTe/iwEx2tt6KGChAUqPLEewIaOQKru
oxlYIW9AvnlOl5D/IM59xl9GmIsxt1elhPlTL6bwQOp0Npkt2d2m0eDg3EISlUIe
N0ZMFbfL8dMnfYRhM0hbr+x9glrdusZf3PvF6c/GcU/HcNp4I4GLU3Jsdg/Vakqc
iaogCChmYSqpAiyfoPgOMaMvh4BuT8ndcbk65xIrAxmeJD0iDE6/XgO6YrxMTvmO
JfFiOnmXt5BitUfFVLCVU8KajLy75MaMwJClGcY7kTZsQAR3S28bAO01EDoboq2u
mkBsjdpf9fXP5V9KkQewCN8ISUTkRAT0aPQSDcFOsAOUHBKFqPKM5cMwdSai7XL7
R4IKmOmL5b8f5Y2xSNwEXVC3KAxKpTVuLP7Vobb6G3sAoYueCdksLKBuhKePmfy7
5CdhWvwCFbCnGzuqaEqHuUb5/T/B7lvlYuOOPdL06HsV7vWiXsajYND/ogHpe0WH
fbsY+iPd1Y1Ql5njNeAYTXGqXzEiih256JMHip1gaeVferX5zhxz3/Kw+23U7SHy
hownPy2NYArIgYtfNK8Ai1e7HgXzDh0q1ZOGmQW2cil8lHxt3k1W/uQrc7AS44ms
QIRSfXQIOF8FqQB9lG/J8KBa4UNE2M/iO0L+ERE4SiZm8QODEIIcm1JjY0yq//qV
f8FTJJKs+yCY2uCi+v/VM2rJK5PQqDDeVBYEg+3uic70iKpFzOmFTBwCCG+kI9Y3
E/ThdMYi72c3BXrErbTjusaEgwYDEU4DyiXZLgg6z1bKvt+cVptZN5KptMHwPuim
e+RgpMh6Q76NF15M2SZJGZkwHUwtEOkjaBaKF5M2UCi3Nu1ph0+eMK8Ow0uQtyO4
c76lZMm3G1LzxYiOuu/PnGtgAAkwmETMpTY5m+r1hsN5Cs21GsR//vQI2sMy57/M
k/lAmaPfEh6eqCyHMapW8iQ/sijsl9FtrD3cQqCsAgw30bWKYkOkIIR6BYRgw9GC
8bLcDAmd9sqPNHbVaQN0NpmzHiMSWbiYyt5CL7d4TCTKM8H3igz7najhz/B2LEkk
/Rj6RnB2vZitOEq8eIo5l8FaRyyaVw0lU5a3uMsfxGxP8x0qzXw1DVQq+IYYSobr
MveA937Ba4zEoevD90eKhgoAvVvzxlVh/KYwKZM+KP062DR+PuXEueL76uXdjKiI
R434zojMC4C6WlCHlYjWZ4OxY91hg4mmydvPncdhsyWZrXRGtt50s0KmRUNNl9pW
lIZ40HaMw1+sJZxQnc7oDVSqImecXU5QtnhXv38LJ6E0qghzENzHAHMZ3HvFSJHI
1e8m63uhhctWsN4UntmGpxL6vqLxBtGxajUT/jNljESDMV2D8MaKRSkaOQMDCK1N
07oXxkH9Vrpu8WedczzuHEVDxr7YYDGFfQSevHuex9i7hDCAb3ZX2PPF0VFLWEF2
TUEmDRCEXvZeN9QlxSyKbTkbValMY90Su40KpuUigTyDJ/Wjf/UageEXj+reXHFx
5sR3pA7eMnLhOMa1+9tQqwZyPgqJ0E+wIjtMyNlMorUtJe5CYVOyi8xOhAYITuDq
NY6FvOtzvrrU2qOSTU0cGkyhwPiSoUhQAzhWEXl8WsySlMy94cpvWzuzrP4kZmbK
aMkpfCoryEbJwRPeuHwyYMiMLijs8JUmcA1rg3gR2Espx05xFOB34V4McEGSNeqa
dbrw5ac0FMSewqjVvPuTKkCKnl1LQDX1YCFT0R+hXVz3UMYJ+UmuR5v6wNxEy5oK
xtcQ0KCkxqUB7V9NeA2k8p9i8QsVv0JK/OZ/RmT2yVyM5IpmaT6wHcKkH+XQjHnx
GUGX0Uv9Bt/l11gnzo7nT+PTQsjP/48qKxcvMDA/Tl1zCNn5ul/PUDlJg3yr5eQJ
qc75zHFbUxZbVhugNmArU1y5nOhFyOSNT+to5LGdz/wW7P5WXqsEXnbsZjNsqavb
z9QpLJE0aefRFVXbKxhxI07ZM1eCFXccH4WIphgH2q2Ecvv7QaxquNGrxZmOaRxT
rbYFFZejIq2k4lgbA10daqqcqQ72GteqikFIRKZMshOC8lc6ZHiYrpMYAq9xSpa0
/ZssRrdSI7jRwT1Hykf/VHZBPpYIhTGYAlDAAB7UXGIuD/PKuDZ7s0wtRgnGzMFu
vtWhw2AO0HqnRu/8g4bzxwB6i+12J8fSXmdUM9kTQi2sUECoN5u+UcOajVYLgIah
02n1lHGx5SjysGlbHNfoSf0EQQfo1yvktGFPw1kMHyw2H78plUlS8VykY8FTpPHO
J4BdGRmB3jtfItXuj6ZUTqygOFSRvYLJckFqmGQoiIEK/PZ9AYjzZaEk9zLWby+N
U4/kes6MTqyoHMc9AD1npmTYOvIQTCjKoDUnpfT9FbM41vNloUDIZGsbKL9VbiKT
dm6mdV+230ofpaekmZpK4M0xyLjSFrB0CGvuJtDmtb3DIAKyQ0iXsP4IcZIl3RGB
aTJ9nq+cmtoO7jN60wb31D6fKixluq15CzSgw3Aq2B89i0x22jjB9FMNvXnjDlDD
wdBcAoyh3PVvn/b9jnKljEbQLOz0Rs3hEDAXAFznjBOlzntUgdXnlBWT4S6Bw1ZM
nYToMqqSoy9Ib/p+1dC2Y750vIwZfgYecgiBAHd5Fu6ILXk/oDPZLnQ1VS9UF06q
bF1BRD4dT/f0WKGghlkxJjgHOFSZ23t8rwx10iVk6bT6oybQQ9ERYTpNYAQo0D70
ukCCZ/jk0CQx0HdgkEIhfB0yYfVxLvzEsBM7mI3Uv5KaTdHFJCLMdm9iO4d095Mv
8FH6WLIhfc/tokMvnovBEMgCelt0TqQOZXr24M2YrAw4hPW+erU27s0e8bxBJZIc
3i3c8Pt47YVZd0MVNL+OtXQIFNFxowu/Aqtltc6g4yxLMP+QHlGX+P9wqnuDbAH7
cqbTCdDVDQCEYJtfxE7EnKXzL2Y+j3QkcMQDjhy+HmTXWprW9WHTJJt6fpvQGTvM
Wsp7WZgYrxxGnXsyp6v4UIkntuOnxWTFYssYs6mPdBM6kNWx6aNfNAbADaDAJc9p
31EYeWfqTS/1d4mw1joz6dAPhHYlMTeIxhySp7vTuYbA9vu+Tk/GGZYc/IKwckgp
rQEtQLbq4OpkWCoMPZ6nmtUGNwtLqKiXUJ7THOOcuGMMDpSG7ULVZUn2xN7LLNiF
4HfbooFX11G2OMniE6T8R6o1cARQ+4POx9LjqUjjitvQZoTufnj7TZ6MCfYXpdOZ
w9mc6uadDeKi+cyRKRBJOEtPlgyaly8E+2hkRkP+g0V1HwZxjWJPY1xnLtmxbA0G
XIQ8U+oOR4JDxS82eLaMOkQTfg/g0Cp5cxVRd71CpFVr9G8ReRdgudLb4bIYBSWj
FFFuocnD6TW+OUr9/WKxzGYAd3hbF1qbXZTVYHnQk+ICM0QyvzPgieaBtDzdbuQJ
cS042jbn0YfG6S+azK2LmPNnA9y5OG7fxyCsA4sQxYfT3Z1Zrc9k5VEolri4j9ha
KmWGGG7ZBAv/T4KnTyK/1xcRllVcFdjUNNTcoAE24kChURRX/RdrqlOCVs8r1T3T
PRKdSO7/hl583dbuc3n90P0AjKqWwWVMKwxZOMekaz1m65+Xq478yOWlWm17hVox
qercorOUtiaf8R9gPqz+T7u3NMfykK4rw0GqduwHRmvV0dXxRdwzn1Q5w7rPaQT3
ryYCAeHDZ2X82W+ywy+BTQGYADVxIWtO+Zhqwa0cybrmHKB/4affye+Wy8Jm1QF6
3oZmOH5Xjb8tQQKHBkmLbNM51Fzp415wfwcpu9G7dBWKOXbfg3bq+x81J0h13ezG
STkzTrxMipNNgFxnvNszE3lNh85gZ73hTuC6NUzqprtpwdt85UCPjQLunA1MfBxO
aoGxdXP8/PfmjDEXZnVz0xLCudCwS37jt+ukgCHUU8apqTsz04CTxLmxx+rJdaFV
f6pzhqfsQbadB79aKnjCvd+KGUTucv0mAT3V2JmFN7kHGuy+jRqaoLoYaUw3lnRL
Y68MCu0VO+TZ3KJ0HVAnu7kyyOdp+nXD8osOZRPY62oxFU2AAlYxe61LXJRTDzTj
C8e34FxTLZ9AS3+k1b+eQEtDZfUs68stXInklnhBHRLyYeLsljwbPYBuV7eIfmoS
85LVmy3WdLrmNEzOUgVRkTXzP7fzVZjmSPO9onxkbA3+NGqv7jd72U6CCbCCrr1E
RGeZvX3qFzS7oyjn0dvyIIUDJFc1lznlVNp0vv0QuFWEyyYoyzZwyMaoonRtpQNh
hRdQ+P9LZDTWhoBJ5CSC9RtFHxwLlp29ylfMMushDoSvcUdRUNEIOUFeg1dqYxCS
y9DOEBgW4YxVnIFCzqUmiaGYCxyoQdTbnZwlOuInqzKyM6+3a2gBVD7qMzdrFBCv
xFAKYu9cPWqC5UzJbOH7OcN+Mz/KoyRD9tjrytIjZ5mJ+l8WxClNR7Qcqnx8dLdM
NNUvUeD+tsc3lN0oCi5BEfM15DnWV9OyBJgype1n/JLD5LRTL0Sw2GLcLqoMUWNv
wnSqF+ryjLLfq5cL/rhjxgzWHkNzS57RrQi3QkC/E3iT18+q0aa38LpJSd4/JXIz
VJyl6Wcqh5tMcCP+pIiK9yesLPeWkaJHVSRwQzZVLPoOXrgd+L2zf+Z4MIunxkx2
7ZKhy66DL1bGNW20w+i4YoRCw/+mxi4RWoShpYwSsFGJoK4JY48uPUMF4CBayNqf
uLhFy8f+k/xYJNb4+jFvXNj0RELW6OZX9M6AfhzvMb539Eg81xqXUjBGfQCp6rga
V0nF+tgIQcv4b7+bkptPJsqus2fbKBABZXSW8aclNNtZL4sNwSlqOLu+SczU5eNq
u4kttBkjNPiasG6LGs/YP7Z9SscdtepHsA8WAVDP2EKdZd9dwWI8jl61VEjujXHr
uhd9NVdBVLzkk35llfdcgav/aL3b70hAGxOOtY34ZX/IXNUHZzutA0g4y8IlXyuK
q6aiempVLaAroEcwzL7dbw1NV7lnyAEWE1e6I2PNGdRvKZje9kzXepSTk0UWa7sb
Za70uC18GW3tOGx2ypgkbHKvhi/IAHwFq9NK7DjwmecXk0lxIj9K+1q34LGoGhDP
59O9pZLdqlRcEbOFDLY4XeM9vA/BmcDZz/4I9pTkAwYJNttnZVUGU1k/R7M5jt4F
aUsorRT7VDYADuOM6/fAuMOn6RWOk8whxStjqYRvqjPSLpM2oHSLjSYssp28oYLf
FOQULDMWRcCDrTtw7OjhucH7SBOCBf6/SPelfBpOHP+GbfHMOpbGnsu3XA55P9EU
byV0LZkmy1xAcn6AeueJvPHmp07P9t1hRuMlWOjZgUKZ3+EbZSC1eBqbCgTodOj2
dUNBDM1YZ4XpLDWepgKq8PiEbvp+7fWZMB042L35gzDuFcJOsYkoTWVdTLtpXMRR
R4SMyqWT7kApuG8siHPrgsBKun6sqJvPKEoc29zZBllY2QlC6uxvPezt1r0CpEQh
9zjYW8d1sJv0HSvGlfrjpqp9tje5L7p4jscuiu4ewVlbALoyXC0qqY59XK1uAcrp
ADZ2gOBsMGYfqK8rpjdvpsyUvI4ODW1twyW2MFzLjXS/dj5o/onONCxy0xy19of1
frj4JfMUhL5pr//Mqh+egsOCuFSUH8yXIgz8UoA0IEd2iwncKW4AnV7yl/kt2n5u
pkUx35fkFe3sfufb6tS2lUj9yZz/Hs/TeBkeC2x0fKBFz3jT+IvX8jzSUfDBlwv0
zw1xHGP84URaYb/RZKGJmMHqx+Fti+Qx3shR2LygdAZhc3D2XHjyNKv9YrBqlS4I
+MBIdwLT0AuCbZJAR8CpLsZjFiSWlL+W0/KED1i194Hr6BKkufi+V0s5b46YwC5u
0nRrHJTk+hjplufvpeI9dqH9Ydeg78xeg/t0EJmMj6ss7l+FxV87I9N/wsOA6beR
DTgYHjqdIx4WIGYBJWnp+kb5jOCxHymVqS/jAuWYacKBDh84RJk39xqK/tlSXs1l
VK9rC8q8dDv7cYUNzJ0VFH+DM8mepm/7/QCsXApRXFOy4f4oqyAkkn9/Q5Acn+Zg
+6q/RtkNN08bLC6YSUOoB15TH/zjvFeNO5fpvanUmEDNj7xTFkzsb2g0JDINoQVQ
m9BoH7cV4BWb0oq03FzXOoVPAhPhD5zH9nieb5Le0R4NGhJbyP5orr13UsMss06l
4hj0NNlxBJII/RVQPG1gy5RR5CjbqDjRY3W42fpAiRzkPEqWadexJqCKl7AFLdi6
vlv4N93JfjJH9tDkPqCC5ojICsx0OOORIDQ27th4QBRJUxcRAX+hcPIy58nwIdMF
e6tDhI5+TcEnnqu6CCktUF9+ReQ/rMx1vW6y9VcYtdqCvoW1aVrtVSSaw8y+Zhrq
OAJqsTb3DcEnNExaguV8sNuwA0ssGMdC+vTOOgGoD+mp/fxPhiTzGR8WnELvdtf4
6g2ETL0MWVimuV5sRz6Ct+3JVfMQQSC7bwpru3IYv6QIsI2QQygu6LCq/2YY7O2D
3Ek9Uao5gO0AJGtIvnv+X0f54by7/sRPrzkBBBIc46/l0OpWyvt2WVNi2hMKOiHv
iWhMgbxgZkWkItFfsNRM/gkx6yzOMnB7ZoMZYA4JtnFlcQEO2HGQZVMfksgl20JI
2Vzk9FaPVrTCjAzPzBq2XnijyqJMttRHo5Q2t5litqIQLiZ+TcjPvKFnGktgxQd1
fAF0M36mbx3ltJfu56M43SDOUKvSf4jeNd4npmdrI6pJqXkAUPKn+g5uXeCgQ3Fm
AFrffmLBBQ/9xG937dJiAu4K0zqLT5rQ4zks1oJXcknjUQFtXpSIdHuaUw4rSF6U
YyXwnAddp1NdCAOwz+4vZ2whc9x2ovqHpze0ANWEwSGgH5Mq/efFn6pqOFqm59J9
skhlnbpQaXmSULjY1U8TDe3RTwWp7eWGUmcl1mNa/Hzc4LVPxu43Sgxb7ZjObY+e
qj7EiUCSzeYUM4h4lx/0aTzzrRA9wsYWnDll/Wt/4zaJFKkg6Q9bf+XshaixLlXL
g8Esu5TaEalur6h3TioNKG0HkEhg29kGzIzmDNYqqnLSklEOKcFrgbijzUlVBWso
hF6ZXEbOoW0EsUtWbX2n8DUrVVMdcJhZaY2D+Fy5OvMDZoNP4SUS2vZzsEklVgq2
9IxPHOwyD+Ng34Kp5uINgWp9ax8dhatVajnPT9ULSSqLJ4yN9NyTuzdBWewp00mb
PnJvVYtZfoetPTlR85C0yThjPQt5GNBriOq6Jqm0iPmpJTRmnvkjvhdAXgrbHPul
eyDHP1sqCIPP0ftqCTrdW/Nky+ak1oSYDw2jEFCk0juDGlpJ+gOqNh8+166RzW5E
ojmX+uf2Fhhfuw/WBioHK1iyuj/NFA6SCYp+aFLv19M4FloAxTTFHh4f8r41kBm7
s1vwqNLwIsEwbmChUTki9ELxhT/WZ2vGSoLMQ+kcH4CJSrPN6vKfoAHQrrqT/zU2
Q/HBwmYIVa+i3wSf+IfpZCEyyGdmn0Z+AvS4puRlvP1v6nfbuTzwJUbwb13tpNWv
cHorE4V3hMCXoTILtKBqwYwrFoN9oF2kQmbIzLT5gU9SCuIseoSIuxIQjf2ePKgb
5ju69MNRB08YUdfGj/CWCT0HC77aqd9nEaQDxOxTubmU3sSb+CteI5i7M8A16x2a
4dtp8C17WORnAhBXABEZYDgAwGp/9z16adql/9qxH5PqOwYxzTN2LT70/PjCBDoQ
+uH+J4DAkmpP/PknDZlFaVK5aLF/L9XWlPS4DQugxJGjKpX7LDJ2diH5NmO0hSzm
/l3mfq9m3kJIW3RXuz8mIXij8OrxO3K9NqOLvDqqkSVuTvr3PSyW0vJopFhiPigD
OQ/xY7hNEBPRqPphK4x7E8A8zelSMp5hndxmrnTZLCHgt28/71Qq7AS1P+HTbhmh
YBaSTWXrTGgu0YxF8/rv4f9vDXRaxGWvv9H3VpjKOZXWhJR4IlDjK+mxi9ygRo0q
zU//ltGTTMoxK7teO2Uef3SuuvLN8y43UBG39toI00uL6XI0ljJi1PdABmVeVAmV
DE68aVnafAiTiLUDvGBQYPi22/Mc08zrvpI+4kSk6RVB51ALACvi0rGb8VKRaomh
0vJ/1L+y3yUlWYOYuuVVKDdpv7ogfyVulEkOod/IWe3JBxetOCcTZERz/d+vaKTd
zxMdjVwIvl2dlgAujXwqAl8Ct60vAebGHSlplgEtURMkWyqxI22G7VslGNYPKTJK
DFrSZSrIEtrNCXezDtfRAbg7nTbkQaM/Gge40/nNxmZoMvezY89+bbv1l893fhUi
sBR+uWeWV3S1qh+JDE9nVvRz0TFc+cyt9KSlBi389r+tUx9o25XDrPeDSsRSPn0J
3Oq3UuZdw8RXB0OlkKZv133WvtyUAwJYfHeCqONP4pEy+N9Uy9pb3hUPK7R6pfPD
2fBwp5FuZzQdZgpQwFxIy83wrlIv5cAFlGdFHLa27kNNl+ggBJ2qsuYzPbOez1s+
OXqzuc1ItBBz4fXi47kuFanxj27VnAsMt8kn2SNw9NgtXNR7LEmarhcd1zZqfpLg
1latoNqSMkmEI9Tg9dEYhjwVa5YtcKvJ8C4WfA12znQoc3CRCiW0nGYbMWp2aK6H
a5ofxKSH0TOAcxYfV1bY6eep2wyOFmYIMX7TsKazJGon2Yb8PJuMs9mhhgOc3n2h
bEefY9miDkKf6YxqCF1LbgXaKlmmNSxA2/d+H0DKepVi7/uKrrBf7r0thGfVxedn
t4ubpwOXvi94gGQzREqoSfD1pmxdATTEAWXd6pwWcHlHsv+4884trX6UuVMcCPBf
9ebmaKj2SwjkxK2GzYIkty+QL3MBM8wxSfgFZdeRCkT9rq+ALEqSkERYO2Btgel5
lBKy1zhYklto/AY0gueHx6ojYyn0p+qhffjiAnvnBP0T4K3yiXJRrJp2gmjzkFR9
UcrRSw14ShbnkA0jiW4SXpn2UslAZW67lGmYS0qdAS7BJyqAvyjrP0cMGHaRT9iV
3SalfNYZ+t3x4sW2XY7enyu17Spjya0PqQezbSWhVFArZMnQC3lROLk0QKXyzLYA
c1Bkev663Rdl6n13ATWA+geTiw5xgjotKLQXNJrc0WJ8PWAqISZin7LoSdTuFTzI
ZMirlikIFN4GqUvQ1nEmL20KWxpwv2gTiCJZq4hniIwdWPBqkajTJuCNGuzCi87c
H9UpYHSTVRt9kwxGgkpH6w0Uqoo8yNLGY7VJ/ESxiVZISE1Tvb/orqEIDz4K5deT
XRh6rtCboWpRm0GmVFAhIzvqsOAfbtTF6atTragEEDaCPhYSX0ZFSxcYIY22w/tE
lx+G6D/RxJatkxgm0+CpOfJHjzSr/js+0O12Q3okrVTra8OtJwwrdWC/sloX4YVZ
IrDRvzpPLlcI+6Hp+WvhkhPngOCXC0AGmaNg7OnjsxaKZQIdpJE1J4y42dMg41wZ
Vqz+lyM+VUoL4jYqBoo7MFnEvqeLvShKt1DON3BJx+LGVhK6TAS5bZ4T1ChwK8jh
oNOGcep9cwLp6SMv+IBHgT3DfaObWrsin+wOny3WwWseJhKdqkeImWCPVMZkuoF5
S3uQ2Ae8O4bCsMppAi66fTM01L4UC5icdppQMBI4q2w1ac0Pk/4Ku4DoEPz8KOIS
ySEsGvshVIAwnKEoQG9/ZQA81bPqkwwLw2tQp+acU1+QSMGTC1RL3UAol7UAQWq7
VOTN8kuMHucbiu5GuPFxLlgIJJKk0LT/FqQtA2aL/xBUpLVpD8GbCRfuK1llQFxq
lMUmeKiIynzKA1kf36AirF8veuUi0FUd5mfCxhXuAomliMCT0s1mx1igUW6FW+0s
SVU/VqbS0EDlZZF70FIXNppWrgfQFas3hxBOgEu4bawhx9U7GrLMJJw4/SpkOGZp
iiWaCaaGfKhKGL5jpT5pKyAHrZm5vzVQ75o8ZUaFwLrr+OL83s8rC9z0XDDbEdJu
1zTZKXOKIUHIARc1aLH01f/pW2YahT3zmJj/h25CQoefyADNsc1DttPsVji+9rVY
zPpXRZ6GS3FQvnvxcq/GVEUbojnrj8yTEnq7+SojaAvUJhQpPWX04QSCFS2fjRbQ
aRdutEq2tyK2cnuexVdJFjUD3VkGatVmnlLjVUj2XqpEAGOmQ9r3E0GuuLICEr6F
V//3E17CAYcHsg//x0mYPfG8YT9Jc496MH39zdnfGuWsB2hsqNl7wJT98NNHbA2n
CYnY0S9WzBXf6lEv/ETRDbOt+jE58MsvkdpGZCEWuqvXyxOn6Pe2i1nOGqMc5R7o
Td3JBB2dmvVlALZytX9hefqETrJBLCyI+YSq76Mx3Kf5LIBtN4RDTYcodoREmJ3j
zkDxAN7rdYIr1r74Kceg1aa0Xvr9qxHo6LvKNsP7y8U1DSRfsNOZeVqRQkrPtBYr
9cszjgj9kCP1HHKgf3zX0hO3EgJ6lg0EOyKredL/9172/rlhlAn6xXUDIMDufOu4
hhqKceP9vDXM3NN2e3y1zbB8MXWAVTIny8nWJU6r8rPd9dy5fs4eZkJ+xTBIpzlQ
JyNwUGHh7sQaVkYSka8PhsJvzYWzzfEwNJbujZZh3SV1ZFWtWMQ+WrgaoyzCSUNB
GFmnwJx7tiUd/S7IjWhPxidnBW/16JXcOm27g7uktS8/YHcdYCCAamB/tBLOxhDw
FEFCRHljX+omDRIFSzaSESlKMibvZDvOdeeMJKiyf9ivQBAju2nVW89naHFyGdTB
0E6/NwfqJwaoF/tKeJ/xikJo9X6yP3bY5GBUTyXHsPn44DpAjgFQqGxSsjvduioo
T9tQDdEicaMMWzWntDcgHqpNggDwAjw3VaT//ct1CdGQ0AeRbiIBH5Mmv7dhWpYH
rQL9vb5t00dEW/77H5HzmxhYqkeU70UoFXyPmGZYMMuPNSTiJwOaLGJjL6OhFwSk
H/UP9QR0k9iakEHW7U4+ozdUTJQqsvudyVTAqpzADpr+29Mf5I6cg9u2T/CG9T9Y
njI2OpZPavlZEwQhxAKDYIBFFot6kEtRohr8b2KH1lk7qS59AL3Bc2rY8xEw9XNZ
si2LFIDy5tAhRT1Wk5SAeiVFyTS0js9R+sKJmCZw35O8ktuaXp+OxiyfLyJ3DMxG
ELurTuKjWJbTblGlHAHmWHYXkCa9jBrW/V1DjOVsk6l5puyF6OLs+uTD5KLWY0Vl
FzUSYreV/zJaWfG8862GXK2R5Tf1LEN9N2M3E3gVK8QXG9sUhVIGTw6upWOOMGiw
Mc5iJl2Ed3d2mlgs/kqUZ9EyW7PEAc+FTNd9DOOqP23IFAZBM5rnlHs7iBPF7kWP
aYwyPPy6kwaJON8GhPgWsAKjlQ4j9kxfOGeOCVUMR3oFUGZoSo55gofmtTwQTiJh
riIkllj3tr4wNrRXGTcpSNUQpbWV1g2b2eYKtpsvs3OczYnajQEx4u1FpCNgS88M
BcwvrPQHAoZiT/kuy3kAXiIlbaT5wULBWaCccz9s4HBzYSrKAIikeeRBvrE5pNuW
otMGgRh36LZZOhAMbvfQK4XBMeecKRDgnzsB6i1kYIGSZJHinbejD/Odsv0YvUVr
/XwCR4VkgQrzTfzgmYh426nJjsONn+pyYL/acVEym0kvkRAKnO2xpHzE1sO+D1Uh
VYk7IIvq+AAiOR4p+uNhJVI0TrHMD26pNUY3+zJPsOvjK9p30nju11Onmg9mMRe3
Noo5hJ5tbx+tkiQrqKMy1Jm50R6Jjd7Q6VLXrhwg4O1G8QsZgblD4w+y5Dtu6QwL
bjZJpn0GeF3j5fZoOpiqbs5WaKPvxKLJsv4kOhFo7jbOGKz8VwleJ/xzpLgJ/aV8
5rBGK6130botzDchQLCw/5L28oLorW4mz59/rR6DfXKm6vuZbrm7OYF+Dm6+fgqo
HnI1e00Ki1aEtZzIcpHb9c0CEoCKWpe0XyNWxjj+BzrFle30HpQQlIoOvKCqLvbJ
mfEl1MG+cxJT/O7b6tp8UchYV1lOpVx3DwLdTYgkn+pTZHDtghoA6siYCvC5IfX3
W04onZu/JVv+8YJ//dr72n9LIKmCGNeMK0OFTvJkiS7sM4fB2kjbNk6O6vTgdgom
bgC28AqQxqsCy0LcQp8W3lIaMhuU34qxxji/lnU4jRM9P//8gOK0qO7sqxfj+z9q
d7mWdF0CSYoYDEfi3ar1wZWIFfj/F7I5q2iBVfLSrA7SfkaiAtxfwzcaBwiFvkTk
zoaQ3ZnPFHUTyqGbVGXMR51yT7tLkVxrNnKWsF4pZkd89/Hj2serOQj5GrQxmoAe
LGEEU7Eg6DV1/+Jfb7bLnZHub6S8RKgbxo6glgQ1xPBgwLAUM47O0DuoWRKVmaAa
bfpKbkCpCQPnY4xRJhYQMzS+WD/BenBa1cUwMnbGtXCGE9+yoLJqFreby7vPb0bB
d9mMkaR27PBLI5lSa9ZHczXRdVjEIPxkwNoJoQhgTox4LofA8KdLBrEPyVAhf7vL
j5FD9h2r9lSPuXfBmcI36mTV0QMAUJsUFoZKr40uE9702F4V09jHlMBS68dmvn59
8gmh2zrh0qbmHJnM4j9k/YdQWa1fTR6Y0EJFKReMd6+V+ugnqZCBYXWtNcCKvBZd
fwsiJRrOgJ5/9cJkkzauBAzVyhDc1T6Uhuh7UXfwm2nGyqiDK6atSR4N1CkMriP4
zmpbLatlrDYBxT2b1Ru7fALJ4isTmCzeFqa6jAYFmXI7ruOPaXQELngv2sFvWfy7
cq9vMyBu5v3TQmjdX5H5AiYibg6f2hA1Myscv4+sDIdE2Fek/ci4RpfHtHk87o49
qqm5AL/FM4vxOEtj624/CHlCMF8EyiG0OcmhCXLbsrG7I4xItINRpXUTyld5BTTw
IvBfY1qVaLFfT2E1jec/3kfDQYI1Eo08rap2WV+121zwiEyFyCnRcehxqIcoTlk4
EHQioKjvT4wXHk6x+EADhiGX3Yds5H2Yz+cE/RfasFdP6QYmu0AmlclB8B0+pt3X
uHmeDeeHMJLfs50XmRUchSvTdcu34n/frMxkGJolroF73zOeKOP1hmudZggBNE97
fEfEMgu0cgimg94WhMAejfrIAoZkbJn4YmWNhSQ5bkoTxXerGSdVSqU+H208os6o
+D9aFe0dGzponoPLk0IfzO4sSTH3GjWtaIZehkIuSWdRCkOsBMjfnvcXHfKh2OjR
y/hz1VNtzJbS5RBNdsJwuYcBEG+exw048dKHzUFRq2bjtWZ815D0w/ym44ARfgfD
PiGAkdYmxQaJkFO2ykUdfWQZkefVC0+oFkmkCJAAqfvOmDN5+A0Ic5aysIoxcjcT
GynO/4Zs3wXKeHlAU2UlZOVFwjMwnBfpAzE6rdqZ+oxTwJ3LLcEMd6WGbsXfmRd5
ZeBq+UOolXr8VIOZsZCO8XfIKVPeDLNpTaxShwEPc6NwoKUv0pjBlvz0D/LCC+rs
yxtJJF4/OpFob5jvtq1bptBjdZBCMyHzVz9jaaJD7btuDfBLuTyYnc0dAY+NBF+D
rcWMp0lrO0W+YMya9bHonQmTeuobLMjr3lCkF86suBjacmHSbK6+guapEMW0SxyY
EDa4g33afRvaEMwaflMq29eOgYZqohRrwb9Cx+F/SipaOd2SG3Kb1iZ4dGCQSa6H
hEdRNRK4GSbPiZtiN7nMjOfNIXYssK679r4fQDiU+9Kr2iYyJW92H4lKUGxZrwYC
NB+TuNKLFp8B9tm6GonOCXdzvLOoQ/2l5YhU0Bq0WfeuQ84FXw9L2VB1T3Ty/NnQ
U381RkBGfpoTSL9BIupyp7+2LMecjCbYfiXUPrnwQMAC0KUk3BlItMRWwD3BZvqc
fylbLh4MQpOCdFpOT26uqCDy1/aw1Q67qItWvtzYBG+JyKhiw543vFffvMweAKIH
H2/WwW31bZnbvpc75BHV2mu1OEzeVFTt0SQu5ei4htTMJxLH+MVCx3GHoi8AlhoG
3AFB67t/qwXE0CzOjXqRs4XSJf9SdAQG43VFUPMAGoUS9vvwzc/v/Ik1GpZ8id+a
z4oPns1ztAo940BSJObx6zaJj6eUv6dDuezJ+Q4ZrsJDuayNXPIPZcWPlkXlgO4/
d3gm37Z9wovM9kHESbFDNpQWAIM7GUas2bbNvpFPEiwFNysozf8/7beBx7626jCJ
OutvB0QU7h3pVc06HMjqJ07XJI9XM12MKT5yCIAvQp9gEzr3M37/sHExgSFKocCs
Yq9XeFRGV19jxstv5/pSgcsYGTqVMT9LjhlUuisvGNFYx7eGSvhmC/1E0wTd/Cey
p6nU3Tf9+s3/zFR7/HCiHNAxkTIzrgE8NDwOeQTqpPYyAlXeyXmQSLfyHRvDBhtC
Xklet+NfU3vfodk5g2RubIvpW375yOhhkWN3vXRM1UcU2wilrxLQhWNPenQNMgo3
nQeEYINb0JQLVhdT0Zp11RX1UA3uodhbBxFqc7HZ8A2BBxkTAqX4bKjSRxrqbkT+
LpYGaHqh6WEgEx8l+dBOq5C3xrF1RM2WHfUVdqZ5tR8/inGqzoFluMDboeta1l0v
gIMy2ZqY3SRdUG1Zt9lbKInT0/fWHPTITX/EaLFiZAzR31xreXROYXmR3vuJqXHu
adNp/9IjBwJSdTsijLrZx7f/TScKp7LxEm9YY7GnBS7IrcukqPD4Mg7Nb3VHnywX
HhevwIhI6B5jTXncIHJmizDbhG+fwmsCjsb3uusOS0QYR7K8Ydyr3ivPejWwe9tY
m8JIlL/s/oxUgZ1LiCSC783RKPyFb3jh2FyBscD/BVEV6N/UcPBLFMDuZQyThhmh
m1TvWOa/H01mFjYAptKaDvKo93BDzS7wEGl64T3kTDijfvxCF/oO/02Xf4E0eSZB
C6IHCC3zr818XFMs4ppNIUJOYaTeto49lnnNRbwll1+fAAuoGLXL/KJoK8HGzZlU
YuG7l6mO0CrzYjaQWcfCtiH6BDQrkoQBGYIaT1PMzea5dWPftYWRh5Vj+h8wTVoJ
LfyW0n2AKclxHXcxbRlRAge2sJ+bNHkc+gF/2E82/fVtADHjcN985l5uFRGhZwGG
eV7OS+HEh2IQzayGxps6sYinUwhU1IKb4EubfAovJm4GjzWn9itjAXTZZCPOfpPZ
OtZyriMo/VH03jdzybDwhhBgpSFfdSPyePB4oUXktvOLB+OzN/Jlx0veiz1Ibsnr
bk4OLABhm0P5+Zxm0yYFowLbhZc/ldrabb1Welm7BUE8ogth49cLho+5I8vCV55P
3MTrw1JssuOQJtE808i8FNLxckgVu1N9MDuMgDNyLQhtv9qaVeus+iXcYrvTyq5o
2lwbVlNIsfUNFJg07Za3drhgP9ulqMY66my0wF73JGu2nd2JQUs9Alyz9EUdA5Ed
PIHU5dmdDt/YiLTTcGD3A4XTa92RfmYbyMjZQBPU1xE5aLGhdFjPbSiywdD6317h
IVUgD8ClCMT1XjVxb0tUCiIFyWeHa8s5FO7qWpfZROw+dpkdNICWmuTZhZ4hLXf1
4ZYqddfa8e6C8mAXCvj3qWP6g24wQ5QFExsrqwj9vQRXp4fATmIwZXjpRZRuzT41
MppMqQm8S561UAMF3lPSAQvVRpwRINaItbX85nGnpkonnZ0DXblFYQli9khbP3NV
dDEcR0qiilMyd3vp2pVylNo/flKQIo/3Lk/cMzmK6c8/cGfyU6MnXzZhNjqEE8g3
7WzJ80AYa3m4MCDt8uAJyaMPbB5h4c1/oAAbRM6ku+Tu9CeQyG+SAGuZTsQ0LMML
wK4BBrKZQiiJ88EOXn0Zv+wm83xap9TqcHQgTVHEgN63vG93VPPdDywXBlt0X41Z
WIRgxK+hd0NF4Ibv+EM+1cVDsXH2SqCKdzvrXYYcmKqqjJQQTGJXYIGt+kBFj5KR
gI08op9xCs67UuuQxhxckM61r7PX9S3ykeJ4QJaJlsolPh7g8e0Vlv83nsWxG4wm
7yKAmWIbbswr4yadRbetg942jth0Pi70TpsLcjEh0iQBL75NrpmQiC6EigSW3cwR
o8k20dL13sMpfh2VMq6D8y+aFamXvO4IrgoyH5HicAAGYmEgAFmTPJHW2gmpYMv8
1t3B1dRmaQCQSxt/mLhdwSWCW79hXmDLzgVo25IJRcMUjGjIDS/8NbZoZ+iyX/O9
VpXeH4lak4AvUHOhl9xDdDkWDhdbKhno8o93P9jqoevTKT9J66f+YgaIsDCulm6p
cox8QP4IX8sZgmHCpo0OZR3riEsh0ehraZJqqdLfTYHxXF7aVpUAI7dB+UY1jqmZ
pbsO4FeuG4K5DXqlCgO/nNZIO8QvFs96FtEoy9mkAngrBAqJg7RYIlNpjQ/8ddpi
Sv+qFc5xWYYg2fwvsD3QX0aTLnYvm342NeFCOHdYGwDKaKnSekzMQ1FpJqIQo3jZ
v3pDmx1HTIypGf8cW2C5Y7z8RklEAP6i45dcFnrJWJeZ/HNv40Tik5IdCCyD3zH8
gXrKhRCpZ7513r/OO4yMZ/+pEab5F9PZL+qbJ15Zl3Kg+24HGmjTwrzv6Q3bf/yv
I9zk6AuTWp2qgAQVzv4SI73vO1SKynw49u6rOLbqCcK9d2bX0G8Mf6l9vb2JCcjn
Qm/AG0R7UwbR7E33L5TLDBI2z6ydsrn8sjx6GI3JX5ksXDKgqHfcCfUtT40hY0dK
otc8JDwuIEdC/mpAEbVxjy+qde+plJb3JGXDnwccjj7XrzmcSoFhD0c18JT467Pe
xFvKIbbZriN9rliL0NBzOBhKqQ7IR3BEcxLCdQOQeK9VkUV7X3nbceaK8TRCn25x
eUE2n/YLFk1hkD7dyDFPREKNsQ//pb6XvJmqpiJJYY4OmKVHtZHhuRBdzqk175j8
Xmcb64sqBbxEvzQLziLdukrISag9IhPCCOYuouoQ5s0qbOSSVbaCSEsLiCAV7Q4o
SvCd3U+JyP2aG7M+IS0NMLO5aOTw6VQchpJLsvPGSYgIX8MHkYu059bLgxNpj1iP
khXVB7UPaAMOBi2HnHM97o/e68Fja/QdYWUHPPTqx94PH0hBIifEDZrK+H5thgQ4
rTqlr7p1hoko5wQwdY+MsCApS/69njll9MIIMMDgUjmc8bQY8G3xIZGsvaLi7p9Z
VWPsBBnkPoygQXGA0gEb5CMfXZX5IO6fb4dFPanNK6vCmS9cAPcLAuZJwiSGZ0Ut
4lEpd4vCg23O4WpWZ6kNAogxaiZDi1PcDsGF0oerhFWMJ++xSPPL6RVT0LY5igcX
mBVN3tIbK8k3o2yxcPusPf32pVzpkG8KgB0SoNqPKIwBNOYhgYluCgUPvkpe62jz
9GefmDafnVTXFJ5YgQdWtaZ7NF5QvxyI1ZZ3+QEiVN+yQku8x2zdLr6829ePE2e7
GqnLgkVD0ygPAROvxnpG7G1Am6lhx4Php1A0WR9lRWYaMe+N/98qcvUsEp3iLXJX
g8+fOQkBlwzhWwNOJtVVqSbDIRQ0MRgD44YvPSg8OHLSEa3BRFFCsc9TD1QRl5hf
eyyIJA5R/2oCtPdr48OXeOVt82Dm4ouBhSvD2P0b/koeMuCAMC9Jwdjaj66/UZYM
1cS4Ru7zZwraVl2I6gLvrEASOewgbbxabAFJTRy4wubAl9x4PFEr1svBz1KtG2DZ
Vh/kIVXkJB7H32rQGg+z+KWMIQmFCM8Nb7mi33nQ38dpjbDqXk3RtXziiZ4qwcJg
UIbhbf8c0nLTxdlDOv2J76S7LnUPlhrA/cmRQhQx8FO6AfDnrMLO7CyKhoS38mA5
qNiX+AUGfWL0WIvsrWVDGunb3XgYjetL6i+fx78+ISYTEKikYbjCjfupbYr8m0Gx
61LCmjk3ZnoueHsQ5hH6Pzna1o7su6B7P8EbmrwUiVjI4OH4edglzO/bnAjevC2D
NFdPNmPicRQQF5aF+FK54UR7LGKOh0mW8ucsoRRo68vl+CWpCzXSPqgIO/X2e4If
03StRcRy97j2OJ6n67CzJd91IraohB3HkDH5MlKGa3fU5al+VawD6cWsYzVwI7rv
8NksBUC3Xmmk5Y20I38WxQPIUWJDpTJIXA2tp5MZ8iZ3I+OHTmoXLkIqqu/4NrOn
VfwZo6lfig2kpzOjxvt2KPakVpLndz+Xla9C6/RC8PGxJjTD7mGv5HfzXH7Ekdra
ElqjiOcPV28bKAF51tsfr33rQHcBm0Ar8Img8Lio0y92aZrJK9dfjgc9NhizY+qV
EFZm2jdZf82gRz5GTEXt2NBipfzzy51wDj6Rty243VYOxpcJ6Y0dL5o590wNelXv
riiuVUNqYyzyqeglDnwafZf/6VHjEjckFmf+5uAfdcKgUo3cLkk56fiKTJ7l5DN2
Nkn62TqLflhuajOvwViXZtGQV0AcTISWiiG4Rk3zogoqmCPKI9XO55bGY7UDezeX
5+MfVUC7b0jNVdB51v5IwBcVk7jMPO54dJoJm7LyKZkPVPt/pWYeayC1FBu5SJPY
3A9ML1jVWaagA1hxax1XlK5xqdaLABNP2byBmLm3EmRgG/qODIlFgO6sxUOxQavK
GSYGKwNzmIkIVlFdLe8pKStG/7X6ATIWNlEFdzreExEO0JziC+gTx1bzJl/mILFP
sGhzP6xhm/ylBoG+XzivjnmJyBzX3bGyTyJ0J2saPN5EbapDKC1Vu09Hb8PzAhBR
Km1P9LCGyS2LeH88R3jZq1QJ5eZFWvFFfWU8EVFDrK9558GaoLa6XAwBe+QMT7Nk
ZEByEoOTilBG/PHAJeDhkMeY4ac5xG1K74PwrpxDaH8jzFSPmKCK9NMMDsdi1yR1
JWtfblcZaxOQSrQmNaZ0tgPGBFxjE4wL/vz/RNxpNtTMIHR4x96njodsBUQAibx8
eXnbJONKWxcnttzcDMDde4Sr501a/Ak2Xbxbdxg+9SbfU033fgep3mxCHEO760PT
TVbWjcIOamzo/25gQJAP3L4aRL8I6bamyRDXOBkHqHJYq44LJf3jix8ShKZKb5Jq
rLOhJHwH3En9n3mKnxt0QIG9P+U0qo5nG+9cdR2/XBPHAaXDEeCTwfg+J3WG/beP
vAZphMVvibQRUlHdrRWCIeF6oH3TFrlBFjh1W9FQ+2U4pfKvUlzcZuIeHaSw0pAV
LimSKNJIyUxm33a3t5KHLI7WMYjaKM66fXuVLFFnVs36QUvIJ00ke36UKKXsYFGT
Rr3kTM0btKMKBZvyxux/tEE+g/mDMPOBtwaIUvV5jqL1VH3Rt994/NeitGJrNVja
mGj0KeKOJ75R1V838iGSrvyfxgyd5+wS8RewBSUtDS2mb4rYVW/kNUnGl4P38FRf
gskE2KttgUAKYgZEiIMYZmr11wJLevRlGKX221PBrvc7vLGNbW5Hx8vdwykLwa7W
CQz14r5Hgg7sv6jbEH+/l0zeUnOlT3KeXyuLV6FbtQcNhn9fFrb7v0+PleqoFYYx
UuaVr1i0Lsxm9vQuUwzd3pPsE1CW+s7fKIyWLSA/RJ/MZfZeHu8oPSI8x4GNwrVq
vqmNNZDjR6bu4s54WBHvjSfafKxQkaol5R/jriTNrxHj20qKg8tj7XARGqU7y+mQ
cQC59NkZzyPNvhj6tnrKxopRhx4K+h8UOOoM3oa36RKD2PpmJqlkujuIQmqZ3vxG
iFCsN4gwkuNtOh1viXILyx359OwLJdOjihGrw9/GxkUzFq02CNMmFDFfJwPfQrju
zCZFSHPx7RIH4S3aoFQFsfPgzujdTR4YZr5aZk5gJE+z78K/YsSQYKvgoW2/bJel
KMyBrC/D35wJxpToFTDFgV7UdjOIlq2hqV61QUGDwLPCdXBpXB7N5UPd9057CNWH
xzetzIWZir2iom6zy6YaVxwJ3Bpr/irz+6fb/P23CFHCNlWUKPzBwFwTt5/mKtPJ
tSrortLMEkrbUsF9ayftVxJgUMbqsfMZTrVuPB9dv545fLa+D0TWZ4013O+7r6G1
zNdkQDKUBB3ZLoTN3f/2onjmM6KZEul8tSBtfNC3Djwc4ZSx/wuJcbxz0M+g1yWS
3M3I4KzAlyRcb9FMm3j2PYIh808OAYtcV4XZLwf4aZYd9BTk+jaZltCD8VHGlgir
3R8silN0aOSxe91M678ofRC9g9Zu9ZtTZmXgnhs9TQW7rJvzvz7LkjZ8AF38JSpt
DX7qnDBK/CENswemu3NKlLoZybAsMnv/v3405vrQ2AFlZzwSqZkSkMiL0x/YrXmY
OXTDx0uMyAr6NhS/iWpB46ZaPR9OWAxhQNnyIZBEkwRwDwUhK4wMMiv47Rcf1pv4
tpun2MUbcuTWTklM85stqU9dLK5Cc0Qb9vuOExEcdYDOYZnVt5tqgbd4gxLvnIke
DMF00VIKXU+UupOKOtfkLsIg8ggT6YUFxqsb4PLHpq+0wUbPVK++FLC+6FojYPEg
NXXamA1itlmI00UsqXmKyR4+vDH+ZBxFqF3sxH5HqBiJcg3AB3olvCMgxefXH38C
4Nc4iAvCk5xFlmgslzF3oCnA9FfHKDZyQhYCczJe4NCz4FCeNB1v9C4zQnBrA/mc
WLQJ33yruBuz1QihKlcy61rYcUQh8AwH2Ipi0cuKbeTahK2dsOATY/XF5v79VKEE
/eJnNyetd2U/03vWXbHeXeB3c7vKAfDGgwYiYkWz/auPw/Fot/UywyV+WCmKxX+a
geZBMebpyLjfc4Eu1VJmjy24sPdS8Mll7cNhb+HqXnuKJQfVOwzF+8kNylmqIgWK
6b70jRRl8h3KCwIE70yjiJVMKiREKnr3EBz4ucuSQDBrYE9BvbXzMBdR8lnGv8pg
FZJbrj20n3psYK2srId61C0fG8LbPn9bp6DiOi5aHMcISCtMB65+O7NlDNWeXH+g
l3+wiXBXNamekN8UQUw6BLu+kprQmcfreI1eK/3Ed/OGU+F18Fv5NmnqZHUgJG9H
4OfORpxDCEquVv51OZWyWuiLG0SeLauJPciN8MCKhKOZlmBCu3oWb8q1k0D+EDuR
1xDzt/HTIsOd9zdbBPClGwAYLMrc8tsN8dlj6ulnYUOlEAouqvZpEAF/GszGwx7+
rqOpS4T4jSiC4/vp2rRrF+5YdyeaWkFAqKUtbWm4WNXDBBiQzMmoFmhCpRXDCWIv
7AlBIssBRPmjT4Qrk4DJVSxefWCohs0JEzXVTjUlvYvCx/njKGYFFm6gjbHZmKbH
K8qf042IHo/mhrz4MLIsnlFJZJoI5g9fipC/TwG5r/Kmp+ecm4tueqVGlj7ujStq
bfwIIFk9WCt88M2nKzfOGL6LW7IUdQsKOPTwUSJldaCYB/TJstb3LOk1GmkClfFU
A74e1gWqLpTIy9Rv8ntE2/CEQK/iyCKAEyQppOyg43ZlczRgWGaWcc8YGEsSH+8L
VyzH5hkWd/N1KGQeLET62Wh4p6wqARw4RTwgAjibNekVbPmVS9/M11wfd0uZ3rf+
iODlt/4WT8ilWoDioBc/Q+OQ/z33Mdf9kxFWSrAmcSzhEiTbiFdGHX9yOj9BmAlA
pbvw2OqPE1LUb6ug1ikDFNAOMFnF6KybsFdTnuSoB/nqUkWIxNg3QDiCeAXTLYs5
fByyMbcVrLZPOMRDfjXh8UHyzv+9mnKfVOCMoSGVshbI+ZhZWn6b+jEDpjU6RbT5
3dZXkXuqmkN6NGNO0g8r9AsdTrA4s7CNDMZCEx8LJj2EpFTRidp8j1AZEEphi5dN
3TDdRZ+5iE64/guYULoKnZtIt0HD9vrGvVlCsTr5Angz/82we2x8CvZsOQoTjj4c
MNC/eUbrKAtH7ZlJsQ7/4S1DGHlE2Kja/EeKTbTqlqKvdmv8HJkxIz5+Nb4gIWIf
Iw1xezF45Cq4kvCS1CYJq+R6nH4q4wLnclRVwQhjUcmnAfzUgsmfUILRv2vdECTB
5sXPzOHu49V/9+aw5DfWdc9G/X60rKedBa4HnV6iP3CJzaobASf3OTwvT8XFqtc7
g7IYZLzG7n9v4eqBdSvqDOuKLO3FBXhVCXKrFOhmEf1Zy4tV2/cLRz2awURjvLNx
bwR1npI4SyXbKwagBzH9KD4KohkfMW0WY7O+ll4zLkZiNwH3vkEb8IjmLZm1XEyJ
XotYhEAEohdTFlB2fpE/DkGbCcemLqsBq36irPivUPmzmqNskQBhMevZlmiEQiyR
PCHp555FYWur4Pd4ivlHBk9LzboGEXjU+SG+ZE3eRtr2W39CRO4dL4RglaLkojSC
+mzoZilprTP8ynHmxsSeCx4CEO7Ksij+T8awlwh/qYRb4c+fvNihgEfa97GqIxfC
7Jd0kerELXvs/CW5AX7VmM+BTcsBpwxHI8EVp06QQfS7h7heUnW9ewI07BOfCY/M
0a8Y70YcO46CocGAcxzKQpwZuGwX7I58b4EivRlfuIJaT7zpsYsM83f+BqIJqut/
OAkkAJcsGl979sH/v3r7yGe2VqMpoBZmxia94hpYJjpYLjEpm9f4eDAhdhDnke+n
HrEdL3d7oXy2HMzEg1QQiE1ZmRzsSpSUh+MxUxQT7QsEuk9pfqH8DkZ9NlMR1ZKR
0PS7FABhST7phHvB8r7frAqeim/ImV2q2RbahJ48k34OECspgmT1owQZuEABrWwt
Bk6yH1fLUiDWklmYSGWxKtOIaAGVYMJ2NJuTv1LYVdskfIpVqq5eqH1P6T1YzKGC
w13awvwFLQ1jv3z/GnUWN/iwavwm21BH5VAELPJTv9DNBZ7BxtgJX51AMQN9uIrQ
/K0vAz1ZjBQ+KsQ9Lh5pFhS1awmju5JE8jh4r8eQw+iSqHXDNBrgBBDH8bHt4T36
CC2EDNvrEbwP0vsA/mqPfTRR8CcsUsMHq300TkACAbMrb+y2Ev346MvxeF3tlubq
igAijlcPZfRbsQlvn0PoFFRKsCYyWICCkhs29RLcap6s+pjH3WCHdnsUaj3gf7Ts
y5Xoq1Xnpnm00maWoQkxsGwagrc5TF2JnmmcChemtNpH91v+ugWJR8+cId93g44M
o1csjipXpSRUZ72DxhHxOTmtjaiofowRQdp1fctb/UCg1oMp/MSVTDyXmn92AWnw
qHNBRrwbX02KJnZFsoTkbV84zvVx6I1uulZnjuYTe1pGhlQ6hzicJitVZ/VjNuBS
oixFKsaNBkdv1A0C6bmPUx3vTwVWlEcqXjJjWcqdiDPCtVvhoGGborTidWnryuI8
hdfR9LX/LN6aokGAHx8YoykUXpw6su6g6eCKQk1tfyw5wDljOLIQ4/8VB+HsHqrb
vaTLCs8xyyjvFFlYSUYKbyJBCCUAHo+QitT/u3ln62qENi6aoF8KlZnEBfSWlFbs
LJNB2RwfQcEr4Gt04m4AvGyG4V/uwRvCdePwdIumZV5hGtx/0yXOT9RH2Wg8Z8hv
V40lPHGRT5QttTRQdDGeBfG5g6CLLQp7EplIqf3GmeYE0U3zuwhFmJqXJtkFUKkk
1TwExQniyGOcd4XOu+NM+NMFFiHErtBWSTVeXbY7NQIZudu6SULWJ9v0ymhxeiES
/OAhK6IIuA2n1D1gWlXakk5wdR9IwBTJzYVnhr0vzr9tqMeKvW3WxxHUwl2KYNB/
xROTPzK1ikNHPmuFLvnZYZ/dsvFoauWnZfZGYvE3mRvikPWBdqXjR6cuXm812jWj
VhIRDgkicsECrcibK1TxdN5IhmNP+2TMWlbRPvlcLmAJQCo4/Xdw7UIns7blxgbV
cYJBaWsYDt+VZMImeWPXuEciba1w7xt9nRzJhZsiEQ/GRXcW4e7Ctm24MLej8uOf
250SrEn0aWsxw4IESdbrSyIm3aNKy2Q0g+aQshzI0bKsgNkM7USeMjaoBiw48yKn
weVIEyPKZ+9kAYwG3nHPVLwopW4AvuwUbfLzX0zG7ktKB2+Eypy/vweG1t92lAuf
Gk3CTSce0oKZkwr07oyj5B4kYAOBIRZJfKVL4zlhyw4Kba8Ej+XIqnngA6jAOVt7
q1/hD3k6YfvD17QXBBDA3y83Lkl5WbV0wH1BTPQ0tmI/W6lFKiuIW5XkVQhQo1qY
pWt+RwjdJEPYAxGnyI8bD1vY+RjRBVbUMF7wi07Rp62SSrul47WLYz+31BABoSDB
RWCDiULJHYJegu+1XAx8AKvnZZhOM0ueyYoMhnyOOw9JRUrJhbkizahqKB5viesz
CDBrGqi5SRJqFWNl1F1N0aWe0TOl4V3UbVBYR9IUMTwIBv+WindGVj47Jc5gGl75
cBf8swLL1mW1mYkuy1PB3d9xVGzZysyF9TcmG17qXpiUH3dMbmWGb9uIq3gc5HN7
RXpE3G9hBZVIRBsQYzUi71Qpq34xMFOvPDV3lU/c+g9evUZnVa3cfAwh5w1wW8/q
GOylouWiKB2cIEFTdJnj39y47VoKMudxYF23RCQJgwZiWwWpE9Vfi8r+8LKwNVWX
8UVU75Vp93EWj8Lpb2RdUc4GOKIshMOM7xXxrgyEZ0f7RNu2/EZSoD3wxyr74Fxr
I10RUUau4wWuuF0Zun2AWrxSx2Xz9F6hw9ghoR12/yvzGMWvjjNllHXZnja7JvGX
E4a2LP5XsrtkQK/MNq1jbiCkl9KkrL/P/9O0C6E/6mvcVXtqvA+214tbl3Si6lIE
Yx7RJO9Zmul3/Id/2ZUb8mEbwfoNJTXrUcn4C2UAFm0KeRX7UsnQm1C/O8blX1yg
v2XGmNu1GYErDnZ5YrQWj73jSEgL2YhHHr9g4E03T70TYJcfvUt3pGjuRXoP3qMQ
pbt+Zdo4JXCOxn+aRtsDmq+E0M6Tl1c8lz0MrjaM5Vm2WIItZAb+UObYRfZWYN94
pjWoH9CSTh/wmd5K/KblzASI8j35oxg2pVB4tDAUMti5Si+CSybMjUEZlhmZxGJy
GpNaC7EwoMisIHZIqKEVRdhCOqSw20NwBPllf1/hAeATKtl7urjINctadFe9lLup
X3BFxqy4LAseBMkbGh6FbEEVyGG7WocF03wl9Fs3NukhHjhyBC0/WVGkLA0T+JkO
PaVreI7Qo7zxS+r8owGjYp14MvCO0vfBv/iXsARCoDYe1k8Drpjno+sbhATaWNcB
lNAppJT/veTOc9Ph7e00l0k15y2s+VDoUIH38Podfl6eLoI3ezkOEx21DjMuwTC8
6Oqgs9VO7hIfxykd5XCnyEKjHl5hPou/M3l9lgXlChria/U1KZZISW82636/0WBy
04u1/r5yXiGwktEpmCazjxu2/9k4PTcr3x+In1Ar+tskyUjhhSTl9pSQByqwGieQ
n1Hs09UMFvRkhxkk0mDKK9F5IWg1ppyCxz/0KdMl109ps7ZjQ0ViaKYR6rSfC9tR
S9ZoOgrub+ilJ+H32ouvyRrYPaGBgLVziuMR1DZghOUOw3BWwFBNpbufrqiRIQdE
OfTZK47qh6v8VCR/PPYbf+bJlpZC0tiSt7DqxGvsOHE5q0YXhtM9CrJrt6iRvSc3
ahC/pQ5QVaw4rx8QzkC/uVRrWozgBuBBN5HTTf9r3dcl0n7BuM4zp/djrZClNaJO
fXsXgnAYnFVyvYO80Bh8tp5l0QVCu3KzVPw+e2T786NRQ/Glexsf+WIR67Ga0dTC
caqqdE1qacQ+gw7+zUPNnwsg8E2bldvtj5SrJnnEaLBPY/fCol9z5eqI0kMmOC7e
rZacsZkO9H+8dOxlx+DWdpJfkJxRhX2c53nVBIZmCVXyKdfgPhH+ieAxKmHv8usn
qrMIXj6XKfyrUPKm541xLriHKpQEd5e8I+dxQUjyyDH3jb/vJpyGX/QPPe6E9lhD
A/AwV/3rVeTPJKlnW5VhorT57m6wEWdkjSxDXCvXUpygmuyDOEDztFNpqs/MsnT5
nWzpaCSWpU8sZv9uQHFFGDyudOo5BTxEc3A52ZP24dawwrRNyBwIW8NWfKGpZH+G
hadpFE9ymo59YQUQk+lmi8v8eoN0JXHv2BgRjTAhL5XOS9/5WpObNQdAETEAHlqB
r+q6Jw+p4LBS1dzlUGKUqeAjlXsEm9eIpu3BG532udV4T3MLK4Y0a+TREMYtHt/t
vIhjhC9kllseS+sFxm7w+qUEGms871FIqYZ5HUIkUxxhS4E/cr+Ywc22p7Oo76J4
CT0wSQzwqB2/TmcMQN6Nrz8u+MBBXiQ8+EJzUAMQEf75MIK3SwyHZXu5hUqi9iZZ
+4f7LGJ99qiQJjcYMiy7ML5AFwkz2805MDpQTWqlzxyOyW29zW9tfIqUX03Mg/1d
aUJXR6xo8WuE8o/fUIE56zfNas1YCSLGUShyNmBLmIQPE3qTXGYDXfBxKmSgw2QN
uXjwJ1dap/bmq2ibHkEsmCGqeHNwFPsRkWEzPuF6dmf1YOm7Wcxgl47ys3IW5vw2
kV7nlck1c6TsUEavcaUlIs/4DNwxN2p09oSXfFvXjCbIFpo4pxLEZ77Y5846vj9W
7yjuvCpjYILa60n4jDhJQRhw2ZDvG3gRcWPduyriptgNRKl9m8k1QMSmRzIDRY/1
JEHrSjwMuAI5NYtM2LZeR8qvzSSEGUC8MZlF0LN2ooSsOaReH6ElsnQmJDQeA1UX
lAfLABUjgaA5+dFPNeFqrQrW9xMf7zf6AGQ7kj5Rxk4RWY0Q+VMl8LaIXcF+rAFn
nvy++6x9qkq7aQ988+oSfP7FEkYhLJfHoT8aPfjTz9x/aPN1225jca4b9lGmXKg/
/Zmh58/y3ErPQ0tehuQCAX32bUrwL3sRxJpPLvHNQznlqMUg15C4hh5bPGC2LQxq
RlIdj/JwywWqYvd26x/YzUEutbmPIPzjZZw4sXiV1YeJccrc3TkAGjWyT1qcMzJX
phUD009hszNhmtK4cUkM0BXUJW4FYYNidS6WUSDjZm6nIrwFU4dJBJukPuKezIde
Dpr8YKUW2j4iaz0UfZUby8VL5uIGao2OnKE85D6PjKqpwDTnUP407zb425nE+X9j
dzFp1iJTCgx4quJOPfDlcwrHzcyWzsQ6benvEyri+k9ye2E/UT6fRH8hyd5aa6Lh
WibM6X47VLIId2GMXWG4Oxdjyp4SBoEHesDgHJilN5DatUyCnnF1xw2eazbhecXo
h7FyOhJrlPAi2v0JKOyWufsVhZsxoWPOCTmX5iNjenE6EmyX1hs3JK3XVUe2tFor
Br1W+fkDi1GAe9YHenFcHI/cQQKv+cZV1MVWmrnJwOLEfw6OGaj5DrdPegMXQuRM
+VFGEz6jI6mXou+jpQBuEHwFdgJPxjPMOOG30FGkI2Nl7tL2sGqhu63Ny7FRVS1X
C9jeYxBh5Wl11HOTTRzM3iQ77Gp5NQ+FPd9WQdV0YjMiOWnOcdfHBW75O+9jcsnk
uYD9ylPIrPQUec6WjCpRGuNBqNVqa/vW+wEJrppSwHurs1jkLku2m6SUdxJPmwPW
VFGT8wJl3AJ9N2JxBqE9sbNj3ijCZ3XhDymyThy3VO+JPA5oXgrrCt2IXzsMR0/E
pHeSKpbEEsQMnyCKIPqaSE8OgDv8RfyxrZ+i5fPxKE3uK6YBpxj3pmI4pfSYFjOw
a0Fsc1tr5sTsW+l5L2b0w7dGMywKQbzuBeXUBElNKqQRXi1Z1kiposlrpNxTH8mL
CdlhWYqmJbRsnO0NGemoTHaBNkvVJzCdCw5OFvLN0LmR5e1/vBSIM0G6ZcT0848/
Zv28G3y+kpKnq4+A6PzbSQWAEOnWkWxUbbeKbTQcZeNocRKtD9+H/lBiJ8PakqGJ
MS3E62V3NIfHvY/TTcFWzvDnTh9+7Yy0djLGM2SmIqnKELyNEaF+4vjw+P88L3pK
2JYxRewLd5ZrO8QEMrZEIiIpJn03xXkpdBZ2DhyzGq9fXMjUc4oRiKDBxNfORctw
TzbsUH/O1FNukAQxvSrQLFM1HKiKA0s87/fYcHFb/gDj5IutZSceF4UJpRpYB49v
DNr2Zq7ts557VRRNrIneb8Kkm1uojE0AdMCHmHq/kiXgJbR0vJzufGGZzcUlQskQ
BI++vlVeRsL8VMESgz19N+8LFztNBip8siFCK+AKOlHhbPMm7wf5NYFnD8Gg8Ie8
fzzU+3nVl/TQZBxjTD9CwQRwNgP2aLj9BqZr4O1qQirnNmAqg5qwyKTJlq08B6h9
RhH8WGmTGREf8PBnmlzDCglvt3BZo/6u+OSu8Mk6VP9tsW3nzDTCep4sByYgX2Vp
FbZm2o3/qR75Zd93ROnGg3oAsruv9Zc4sjoq5aGap7qzIeJWej4Tm66XB7xZQN0O
RLt/Hqe9N5aHrHOK4c7s+RYJ4REy++uCCNv8vfeMDWFioATFZevjmHCBc6SJqlQi
96z2tuuBRsTyBy5pA6X6RirI/gP5NXwhGEXwS4MoUU1JNcOFQe05F4xmt318k3gb
pNKIvf6R79tr4YaVPMcOB+G0k4LjAygSNubM2uaTGTrv6EbayWXbi/XeifJAHWUG
AYMjfnmPu9HOxqA3i+UDanSFYxsIuwW6zX24NouXI9ECbBfZSohK+PMxg+0naACu
7ixZp+vmUJnB0XGXOfEzAd3KJqWVDcAY+wWieZQzlileJJwoAtL0J0ynf1ddPoGc
ZjxctqHG7kewBTWqjiws18Nx4yuwjrtkHqqTp8rxk8MpwTnFqT4cWxb0zquvIc+D
bbSSrlR1Hb+RfgYrQq0EBP9b1TR8ylvuALdsf6CzLKejmYnaDppQOIBZ8lghUZdD
1jMjMbztfMgnA1eEmNzRBUt9eVIPLy3exVbOGKSZROgzZEs3uvvUMXd80V0sH/gC
27ZheFv3ZiSPP5736yfT+YBcmwoI6Gz+ApTizSiYdaSiT8qc2U/91TYPj6j2cJbh
Ee1MmI1/c5eOCi/MRxO/VsnbtYt88DcVwa7984tDdRCOgOV7p83k48rnjvGys4Jp
rcnHvWD32CAKp3CGhVFvmz9ZW/pUK1SHzzPjMHFbxuO5Mtix3DurDSQIOyaonb/B
BoAr7GvH3w3fptFYimKb8tEO/S13hqQr9+gjJ8coBRugnAV3Mx+ji9XeA+OIOffV
pJT0HE6mciIP9/dt0D/Oddhc7gA+iWntZAlQjvHCETG0dQWXHSOmPiu1eK5CdZJ/
8HOC3ruMA0YGZrtb9g4ONFBipwwPkj1pn1+TfvHVsLfD7wuMK5yQFK8DueHAKO3D
HbeZnNxRBO0tytwD0sFG2/QI+WZHKYSv96E8fKjHwecJIJOO7AZ8OY1IWY7cDrbh
MYfPHu8W75F8hJzfa9mjsfJls1P8lpiXiy8TRl9L7d268XBuLN77NxQLmcGed3nV
nVwnodfMeoRnkjVEK0T8A9V3BLnOzOI719Cki/9eep3KHx6nTPpon8+mL+eJerkN
wj9TR/7+QA3ECladnUVAWt5PXUPsDv7TYbl/5XZRfLuLAuUDl84ERm9DLGFWqyKC
Ir8O1GM+G/xerC8EKFi5M6yv9pzVUXNQdUoTuBxWxuRafrAUcNCfhZCnJS8iZl2s
ofjtQIpMxvwdo1jbBEnwg/dXeNWybr9AbqMyKY8gtRAr0QoWpf9M7yuyq9LJU8kP
wfyu+EXPxOtvg2X1XadfuHxC4SFD9CKDPeeuCQuVOpeHVmRuJhcSznbdyHlc+6TK
YAjw4BU/qZj0EnzIU8Au90GuBHvNl+AKGm6tn1ounJcQDw0TlzPm08aAJHeuR8HD
YvSH+tlBrvSdcB432IHGz4SZBTL7yRGIgGaxXsJgZT4Kh47y9NV77Mjkq2SXEWav
cEaU9ZIG9LEhMHTuePJN4u1TWM1QxX/O0GhJuZED6kX3aBaPYAlqPBQLlvOMqGFQ
Gb2NucE7WgIib9MeD4RrwAHHYt2OCSCLuU6YZ8/VbwIxu/Pu78viP7jPAmTgVXfM
VRrQROMbaOyvn7zu16LKXraKmhAnEhq6aKEJHZZOYEDSfpAf2YoW5o9Cy5lWjL8u
G1zBQb3MaAAsIMKISh6Te1giXQw6NageboqcdfB/OO2sQ0ZYYsV38uxhBu0rqDo/
yRPZIl5sLoOvviPa5RznJ7HJ8SCOgsl92Aa06yBvR02cNdeO4dQ/1aVfa8WQj4WZ
RlsxUb9WDWt25OsqNyg7C+yZBITRqYzvRSpYCGfhSUzWgmzmmyYMB1ELhNpaNp3b
pmWQ9BZHDG1sve2ajJ2m+ULBrHnMzrW8e/HNaNK9rJKo3KwSVFbwQykQb4/lAPn5
FVJUn8F6bA6Jv5n/j4pm34Ib3L/x3sg1zx+NYfOZAWBDglh8gc//oO2Pw58O02GO
D6JJ+FE4xO/ZCKxIKrIWG2YySccOyIYds8lRE3ZSG022ifgIavALvP/IMkiE1ay0
My19/6Jp0H2mgxsKmiTcx+GByrfbZPYwPlgDV1PtO3gt8PUg26zaV4ZgkKhLhucX
40yNIgy/Z5Xxrnp+rIrf/iMzXJfzbbMVOFHRBLIpBk3QyZso/gUl/rmX7DjHGhGZ
/NBfH6x5f6wX2uLI51b8VATk/tawrcL7wJx1VJFR2L59Uc27sP7WLt8MRUctQ+PE
BVXCbrwC+so1O4F1aQCK5sNMCk7/L6XQamAch5gah+36f9UxGY3f4r4GpsR4b/BB
DtRDoTCncjc9gQXZ1qQf3i+UsNN+XlPUDWCroU7MgB0JJap/eI3l+c3ZsArooZCx
yxhTwLzE7KTkpqekY/IjsNiKYi679u9FRuCJg/I2fG0RENWeoJ8pHt0eNNW+2UYQ
ufS9OC+x8xhIdx0cWkMre8JP+XQcP+i/HPyKNaxNjOrqW0xaueDSKJHS80hvq1Vv
vA0EOhnOyU4kBKAgZYomD0Du+gagMif1bi+aJOXzun+F9VQl4XVRdecDWNcuzV6g
yPxQyw9y92D71RbPOn2sHA0FemfpKwjjn2ov4ynYd+UtQARfpMtBkmy1vY+eDnmB
ci/LmrXznNR5qql4Ujdve0yi2HrBGX4ifUj139tZuFm8RRgDcAjyfjCPge6qkVzx
SHTEJeLJ82462v8V324uGzBQfalDqkM0DvkYKfUA3vaqWXZcyzhOTbWOZPEuyG8h
SxRDXbtQilrcP/xSa/rSPBbPoGJrVJykzx3bh42EJ1Z6gAdhspAXezjDDqiNBsrg
e27X9cIn8H3DyKvlvGjaL29avOBGy1/M4/XNdWPuTg/mkWkX9FKA4ki1Qq9YTjiT
k+Ahs7gZT+DE4K9idNJpvqdE2uEikWfnx0N4XWjquLrToSmSDkrOJ8jLtT5xctTQ
gUO1c6u372HE4EotSAuHuF1kJqo/PJ9jcg2WcCDwyL/I25nyRteZp4LZ2NWa/+tg
5GMDM1MTbQGs/L0woDIkN8L59CikYf+MZuqh7pugMiQRMZprbgAa/x50Tht7OzeT
M+urT+l51S/QCIrRxwvpGWUqq+N8ND/BBf7Few9gNujt3jI+P5ojqak8xozgngAC
jX/DO1M8fhuxOfCFbnAqDJ8qO0jJmv+4iDTsdvZaoK7pr42LyM/SbM6M2g0VEvnU
uTT09RE1J/vqcfsC3EFmrk4OzDgrpGK/rqO8h60Ghkv2qkyFkGqDc9oqb0TclCp3
rXT1OJ0xpQfmGfVCJNAsvA+4kTLufD+yGIW9UaFed/LoMgg5T+Cw94lneDmNwF+G
8NFiwVpCFEvCaVnCeIRhyp0r9Smrn8nN/BxJlAmWFWqxwBRmsNvYrUEC6B4shxXl
/lSbfRxIaMMuXzsslNUulTfhAuw6yKscoxtXD/K6JEJdw28HYu2qR5Rywjtl1Bwf
nr2s5onnG22V7YPeQYWHT1FCL5IqGJsSof8VPfXHIZaN3a9+7oqNKmg/yUlmXUUq
+ncjwn7P0/xMkvQcCljKLYY9Xb8JYlzZjoo6Oa6nvL1zVDGN+Dwzuv/t9R/IndZo
u4ammWmDAWzKHXVssVwqCeKWW14sOIYBgYB+WoM3orxHbtBDRmaWHpiF5cRiuzCT
1Cbv3rxpCQ8hc3Fk7zMnVtYyT4zVwMkh5rC/g2L+KxJmCEh4Fs5EPuD9fpUcZXJ2
GZtdt1e2OQIP7gQtw3i/O9xu/yOE4cF4nNie1sCIrrkGzec9hMiQZ9jfK2r8Jdz7
KN6HOM3YdLj4AhanacBPBEGEPHnxUJgyRprXMG/2IIc4O2wB4efIx1HxAS9KWxxp
mI5ELHMnVvRfWRhYlzXk1Lj6FtPBBdK6Pz7DHNGCTqbesCQ4kZRZzJnb+/Ewmaz3
REUJHhWT9HBt+9znIFaI6z3BOCeAnc6xKuBmZPtLuPHGW2bcoafat0/wivyBFN5r
3xX/h8ktfyNDFY3hIviFdwT9UrOTPOz7+I69dq5tHe2FEY6sgHX3gy6K4Fs1gPq6
FGhKuouMqZZFQUA7ex5DaeZYw9kEdMklCDIcN/rGbd4joiXH4FEfezHaL3KBWEAG
bJleCSKj2LSNT7Zto6TcAnUYapkhwSXwHLbfgYuUlV5BGfCsWk3jjy8EhtdZW8le
1b5rKtdjfcXOfE2+TvqTtUzyVl7opTz7Hq2hU8hNkUJDi82lT4wX+VTeWjqQ2KzB
A36vv+Dm65tFQap6XTWriyf291DpLCFXUZEaiPHCYD2VVLisdJe84PV5TUmctBIv
Hx/8dMEbDL1cLPj/EQhMK3bffmXqbxirQMJmzzSFYiegf7reyEuFsMAQzHmKh7Ny
QfWYpxXI4iwMY1rUFQ3XcIQVR0OiewtsknicRTa91Zv7+nbDZiAVTLG2b2x1n82s
Go36LXUwwsR6mMfa8mMUstv336VXgqohFXC/puIJGGayF0TgkR/puzJmkxV1q0Pj
zkgtzcBQu7907YuIwZYNCtghY46gVUKl+dxmJR7rKH0EYg682TGZr5GKkuVLSSUl
jnIscURo2FQnC9MFagfHQw2T6XPHTkhRgP8684MJ+/ioB+GRJRmfj9c9Kl+Rtlhl
UmIx2ikB8aTvNXmQoQkgAIQmMscZ9i0w97bcTqrpf/wb9KXCvd1zVuBQNB1YQx9m
Io9QaC2/0f7j7ne4IOp4VKL3fSgGol13Z2fWOBBiqLRrsTdVZ+CDpJPKBSrla6pF
QGc1GgN20ebTCM1cA39F9mflxFM85FoT/5t/NcGltW8A/Cuj29nWoAyZ8EsswcMG
e5Gvuljzonphhnocla5H6h/6l4jwhLAFcuGkqZyvlg5r7ZEZGpxrjFGy7PDOLFAV
UAbM2mnAISJ8bnYc/nyjIfGsnEQjVXH2inChum4mOouClEVDfs4k0AkHr7FiPi40
5/YZMNayBMu2mvcw7pSPH3po2f94Z5RdaqcnhehsufkNnoIb4ZguKhg+CRuMg1uH
1D7oPc1h8SAdPFobrRlDWnTib/yapJOwFI4N1WUVUSvxDYkIHuU/6vvWdWJDDRSD
7i6jA5jFLx6BRGZtcRv6V9JUP60ZrXjg5ZduA99GGJGmLz+EiHyNoga4pgYPjWPB
pv8UQ6e/xOlC0Y9j53HEZkstrlDsWOkVkGKc6gu83Y2BYFSCyNGwsizByhd5fUU7
PoDLj2PtG9yl5yjm5P8HuqbtIYJhmwoW8yO4AFqcescUFNQnrcEMhi9hYBupB1dg
dIdeAZuzVqZB7OfKqmkVJlfeOb65pNUSLeEuDB5LYC5pOsteku3l2c/J+54X4MVl
gszvORvX+pZkX4xFeBZU+pRhd8YXE/2j5rSSkGB5kMO7wDn5EfoiNda1KxmecQWF
gBCcgM2ekpItnPFwAyg45wTdqxoJUFoYUwU+ZAwlCAZSjky5OEX+pCxYft0428kV
QkBOqR3II9sC+HuHFHygeXV/TPFib8o0F6enu+Uk8rUFih74BPfFRnCEn/ND/mgK
uqLPc1YFUr1TxglGJmHwrUZdoksqZ1G1oaJXzCa0WVQsfOA5ykKEVYiTpu+iNAu/
KqSxQV/igF5K69AaesZBgFSLTOzi2Hbb0Dlaxj5ufp+ntOOkaqTS648EI9ihjVxJ
NIklC/RgTmhnzhE/mtavCjVQVmWPSLcb5qf6c6De/iE/s4goVDPGiya7hiXePFf/
940PA4xJWN+7jb4sfaahJ56mkHc0Xz9nVbP0dfVfOHHxXDbDMavKk4Rs0CIfSHQh
hVHcfnlk5swyWD3q5o0+1sL/5U03JxWdPM7yhVC9H8EWdI590jQtJl9LPtTRXF5n
tPI4V/ZjGEl1Pu7A0cVR0ZXOncKhqP5Z32+jBFRPr3r/5AFHNdmEhjLD629xm2yo
GetRGFR1RVNuxKdfahx+1iIvFP3qFV3ighL4s27AOs/L0URvS2PIuBnZJufSKxMS
4sOenvWxeUfbXjt1MNH6qw+XBFCU9HT5cj0NuQPoMvCJnMWEYTsPJd3jX4U0dd3d
T8NGYwxn+S4EurcUem1PX+qGaw4eAt6a/+4RTlBPLhgCjL41SEiH6Z6flTB4ji8G
ap+XU9xO3Fwg81I/1iwm4AUF7xTr/S8xipZzx5Il6FDu+RMrnGh/zk/EmxSu/tLh
NAXSGgjAJn9Ncujif5TBNlsWnM9iU9mYvbe004T+/oA3p96vz++yQC77TiAYqCv3
u4uWbseeHEmJ5OhtpCSKNYvUjXFDNQF000TzugSLcGpX7C1hDFRcZRY+KDZkX61R
pMHIw+Hm9Xfnv8Es/11WCZO8eaN371RdWi4bUBHKqDA77r/EKNXZMeDgOE6QqH0h
b8H2yLe4W5dnB6hMFtIret1wGx/W2VkTlCN5iwCQoBD8BPIJXMS7ycfvYGAhQWH/
VUNXKNxV4LaZgJozPX1k1T7qRobfbXN57IZkdfJ1+IFM017oYkDgsQftQF6w8G61
NSiesvmS0zLLI7+6QGWWrVcggZbJqWQe9ceDQJ2MuEDyNYXXx+q8qKFj8xeIw5IO
vZnxev4aN6SEnSOBziSZhybZnf1lSE9akF6s5FUgD73i5d7e3DYyumNZKPXZjAc+
JpUljBzcVzKEFRTZ83VuOTw9zzh1ZMgRmay1MvJYEUjmPopuSElCiWdpwao0ES6m
4uo5UZxiS9Dce7AXXmtTpcPD6jvC1b30G+R7ZQkMnCvJl7+6T055S+Io+oVJQtcC
4U/T+0laSf7Qe+w5ug10TwtFqGcxs4UIAbWFltf1JxAde5falG9eGJIolHu6i3z+
zKnstDsNFlBcLj0ZW7RKiA4svR1Ih3tKPOD53QyxzvLq5xjPYWn1wKmS9Xa/+/5Z
wohXYdL+3tXSSMb4TTW1guJAPot8nmZIcHGt4hVrFBpb+9NmTW59FJb2te3OSm0+
Ctq5XrnjD42GKQxsR8yVLoCNxLdHDh6YZfVXqIU+GkdJCGHQ24np9+t/O2hucj26
5bVagLUWiOWtRg6UPXa/J0MLoDEIjVfkYrGY6RyGIue2+7XS8hFhL5aThMFkPpTT
JBKoOIbgiWWlwNvj+3DkOeJqX/t+TVrjoQVarTvGAy1lQgx85JDVL5nA9Jb0RX7Y
TDE69Bh+zxeq3NvPKOT3xreZ9KxeVXyQSCK16rJLgxCBeWb5Hui+uYaZkbh9dIer
WCAiJa+pYz7i6HV2lDr4t7m0varVSsYAhLzMVEuucx88weD0OGVALaQMAaIHMUzs
HsA9X2GVFm5I3ydAq9RvtCjbb6pq/UE54T/+dOsqOnM=
`pragma protect end_protected
