// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:26:02 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AFE3o/N2yKxF47exZe79CQEARUdmFdcWI3uGNcLX+yhE9GTQ6s2Ey4kbCn8r+dkj
BIFhpOF6nabko5tkYG4jVJqwTfBS2E54a2Z61KcU7gAbfXs+7glDnfpePPUWzwzN
3SdHfEDgOlGdTSwi2fG3jqxfoQBDCF10t+zm76Fz4Sg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25200)
NlkzC4cjHUCjmce6FlEUkYdiNh42xf70MXlZtb/UNgaVwzx5v/1XiGy447BMCqCp
xXhZupUsyk402h70GgkDQAs5bS+QC+FfcLvH9umCYuvnbkwPpetnI8Z2L+H73yA1
DCEJkFtxQP/QEyhqrk2OIRVoIWfxHJ/74GU5j6Cu6df94hmneCPqiHZ9TjIjMs/w
uUxCirYcQTNUOqnQ+3yF4YCx+2oOix7n6afc0N4cOYgIh1U0jJCN+SM1odUN9uo5
1jiglttMZgcbOlgZ6juf5NQNJigBL5VMEpc3Wuy7ZRRP3OcUW7j74Ss3sliwLZsN
axbXsEO1ck/GRbrgbFCam36xDkxeyESeEvVNXnp4M5qyUFCe1AuiMeTy+q3xF21S
K73rdb1gS5dkpPtFYk9PYlfZ5hpjJ4WSmRelR+y1Hi4dUoekA6pfZXUkxC3/1HMF
AvpGneU9rKygayYeAnvgSNuduoy1e/Jax2HImOw6bDwkckAOaJrkc5ARytS4zcf8
9uWkgTEQsEONS2vKNoKsGUBdffsPHhUNMx+FhFmXKBiFDMqIP6JjCNP4h1czNFK6
xtBTR6G1tfeTixG/h4whXwJpwmh6y0CM70tu84jTAv1ZcBSEPnyxYpJOCCSLBqes
9VTz/DjQY3HITkwCZ8f6u3ChfG6A3zVVmTT3OnDNNq9uJ0Z/Lxf1eBYhe8Rt3PGZ
2u2UDd3yCGShXoRxSS5KGbkwFm6t+xB7QKeMkISbFEcyNI8xxuYLYHSy35c5UWKn
LkPuBiW+QR2ZRL80StrSFD9lqJ7jxR7nlyGkHMZLpwxQcmOF7gR6zt2/k6VOi6wG
nUFghZj8hJMVM+Gf5KUemhMV6miHon6r24HQWbxoCJxyXq+G0yVoop1FvzU/U9TR
OnVlpEWnTyPZjw5pv7U7reZnAHxTWqEwxQF6ckht9lgvAwBdQBebvA1grLFfOpv+
+jx4l41qrxS1qbCfgGwq4ZE1dwKpV55OkNl+AVe1RzU/ZTskFiAK6RhOPSKEPALh
fH4ld7lZgfxHITz1CIcA+s+AOr13/7Y/BiV/Y3uBh2r+cYALKPvFVooJNGsIKSZY
SmZ2o34Fn5DFg8WfOHzl6kGNSRCA25ACENsuLCbYyxVzb2QMYCRRiy+Iffgfv/xU
jRiwEDLfTNrc8Yt9FxB+3nVTm53gnoRMVcNpQRu5leGGFM7Ql3iIjqcdM871Gn3f
tW6CNWAGlEU21mIEzEo7PDdUqIP/Mi1FZisimqQKbzSclZodjzRXrbdl+stDmJF/
Uh26EoQjTnupk+bSWxPnSEc//t27KXa6MdWn/mmXVVXq089gQ6zJbkpCwZHd2CW6
TCh/0LD/QMDIP7yHQ7tajVzC2wxulK2DwU8y72gTYJSep3MKdoYirw1MNv1oE3na
qtzsNAf3JI8s4kzXgYTZiPnd/Lp93IL0zqMBt7OoDLEkRaX/xqcos3fCBzigmy3r
MJZTgRkRCAZAb+7qSFWy91+Ndk7yiGFTfLeKgUG74Sr4/ouOlh1OXNx7tf2Siqg9
mk6VMWD/Duy1jrhMq3uM9QM/+YbFCMpQH7SFO75LoNH83Di1f6hiAwd6IAIcJAeW
exP7PUubjbtqBkomrQlWI4nJUzPzcgL41diup10ykP+sgGdEEglJKTCcrQ2tQZIO
2eMf9rOJC4mHWlVrztqHkOQRWbkCAFNT/Hm8TyondsRkWSYE0bNT5T7jFczXBGyx
aLJBjmCsoSP26BEiQagPUV5iwtuHRxyjeU75bp15RhzFVEeV+IiKwUR6YuTjtBUr
mY7RegWkD10suYoEk8ATXBBFa9OVxK5V1d1vLsjcI+rvpa5H7ogBhcXoAfME9u7m
mqho6/qz9t/f7UlYVhLqJzlrZXlx3knQnNsMyUko9yUI7K92rueojKcR6ftvfs2L
26aL7jZBKghXtqaFPcpon7vrvzIGi1SYxUySlqhwgA3bjFtg/Mam6M+e+Lx8Bcjh
lZSWM1eq8Pz05jNQF4+6Ka+ZQtT3JHqWOrICb7c80xL4zdDhfMdby8ZYE+iWwnPU
TVepyQzd6VxENFrfvFy37mz8bqI8oVymmelve+QtLuKvYbVo+h7gE9Q/Y0wvW/+z
ZHacFoQnNH2LQ5LJJFhO6kHs/TYRUVRW4oKONcgmvSLTHC7RA56F+MI8B95tR2QN
mpMebq7G5gsNQ1hXXmnyyuPpX4p5qB+Kou1J3X3iWr/XeCwQs5+V6he4HLP/05tQ
TeNfmc5cItBd9vaQxE70lLQqweqzDnMkvCJJncZp+RKM1fW3mE8k25nqsY68PN+8
VQc++RosyxfhtbnXG4YKirK0mxQdh41AqsfhBSE9pbM+/of8uo5C40ONXffKBpz7
iy+76LxTzR8h2VhqwR7xuhui2onOX58Pt9N+TON+ldRiTk/6UB0LxyETsttRpmEo
u9884biyUX6zfLQuAkwFnr6mbdAKaqaBiw5GU/n08hIytnElOzGNDD2QlMAYlgYv
HPvqYg7myd7XMqqmho8jv+17+zUa+0CVN3Xt529PMiuNOEV68PDbcokgMjZD3Gfb
4rCTgfIHIL/eBV8SfSpOcDv6es/n/HVzmnctycUGt/xRsLkP6c1N9cDrLMQe+ni/
deccpvhyMokal3VG957bOqeAMKjAmJgFEJpvR9VAF8OMt4/F0q9Dgmv5eWqQySQA
Xh0zUWUe7F/hytcmZ6mJH+ZBde3UIjbUwS0FubB6C+p397jv1WmJ+YyhkGgB2BTH
CNT6eAHklw/RmimPQgFedseLU9/X9l78qQ4RZuPbs8XPhGHrPg7tRTpyWi2DJxpT
naBt9j5nTFobqlgjYXedGv306lq4F5OingvP8lutR0KH0AhE+9HlABxNlVN1G4LG
CaDTALQ6ywaTB7XU6Rs2rsnyAacyyyG3ZLBW7KNr/DKQMgzfHmvZhuSvhhmYjKGF
xMJ3UlOz7fmtgs1K6rH708Vm2gc4plGqx/3gbruXHfiVvJKjqHH9Jh8fJgOH9v83
43q2X260uOKIMZa2Ybcm24KjdjXh8nYnXIF8HOQ/DNlS6rtXuckX5fsXjIfX1u2N
dgRU6bhFys891d9XKyoSUn0NSn63gfscb8F0xR/Mqn3Xe/WJY8EwDHkEvoakFT+6
rwaMjdMHu1dSD9W2ztPVtCC18cmhlx/nZ0t3gwTCleUaN8IpoPfHJO+FEiTqO1vi
DDHzk8oPQt28Xokprb7AqkMhAIy/AB5gbWSFhwgpQA7ClCaVo0XNODm+yc4wHwId
DxWbuwgAV+rwQKhyxRfMOUDxldYzzxHw/1UhTWtCXHXWnzvpQJkbPe1cRMdxxvjZ
V23alJZdXeRIEhkOI4vT7d8ZfIymKqbjL9BarEkldPEvV+cUUJhlCMmPZ3P9pWUe
l1PhnBNv7BFwIa9/gDm3MJJTRvXR4TjxJ2OrOQiP+5Tbi0Cp3FaXnKfsoXqPaGTL
2rsgZvHULLZ2Fy0OyxlGJ2VWw85Qxcyz/MtR+4vE5PGBo2OVrOFnKUjhDzJS+7AP
rjGtzeixMU+dQd6RXewr9LtW+GW0ghaeNfhXDHCStavme3HkNj1Dn0UEIZyPA1Bb
kdxw77l527QW9Tkp85n1ZRRhzUFrq/ZZq1g14WZhK82nf0RwUpvSRXU2eiIgmK/R
rTy9eHEHnn332EGdYw1c6ajZnluSlcvkH9RbAx5mHggi/GcZ9LuKbIDp8jEM0f/i
jxmWKBYgPKKJVv7WToQhoeIoupXa2JUcV7BFsFrcfAwqI124b+vEpGsAN6SjFY6j
qNB1b/gldUkRfOKuDcJWlyUEragzALOVKkwFK4uVygX7hQN+I/Gmgg0FxIT4tfbu
EMO/Mw9EP/Qq8PyL0td2wVCXD9iYMBtIUD71Idp6XPxMkfj5gjavAjQK0NEXt0Bp
MhA3NmW7XgyBRyrp08tUG2jvxr42GdgIi5jkQ2e1Tm4+e/p5cWKRXxj24x6leqpF
LzJY62ItLSVQGyAq4Z+2zsV2mUYcIfWHZbZIn93g87zXJ2KI4hcBNgtHgtXVwvRZ
xTnGj91av67njDf9GOdelpa2UhoPu/84eLQx8RSZ8AE0fOQ8P2mAdbBTFkST7lrB
QPDgw4CceDFmkFm06cL/SpCux5S66ejiFNC+w8Ph/xU4gwmiX+gRL8jE0cVmv4Xw
cO83UKQsQJUk6AMzHb0yT0PjwUNkXx8g7sdDAYNpnRr/7waMBcPYH6qoYhcknPfW
lghnpx+2S2iefus9TGwrebe0Xw6rkA16e9e920PLPlBiVpTfE2IEaMZcUYo64+AK
3OJyvJ4Ok8FuoGlKhRyjltJxG7GYJWFzxPOo1mXeljHpIix/s1mq9TS392MTFWBZ
2EaFD0cG9aNekKutaJZ8boZQi+hqKsHK7vuxfgyLAGy79iPLyQQLvoBsKe7fPvM7
WwZ/vN9pEug/vFPtDGUMAxtuC/Nhb0ZcIyAqvDFl6lTu3u0/jPJphi7ETX/YtgPU
mbAQPHvqqYGptLh4wZxbCRAvRCHU/WEG9dBY1uU8fSJlwtW1Vcig4f8UJJsKz2qt
MHVfdgPX5yex21MRdkwzgCroyt6HvjpFRZ7Uf9gMqGq46Os1vxjMfjWCUKgNMeYt
7aue1fnRISTQRBwtzgeAHmGMjnzRsnAGiZn92MXzAFDQk0vB2fdOBIX5SYPq5QcA
fAMHMmQxSf7vaS7glWzIqPVusVApLH/K4MG2PuoMDRAjkSnxDC1XNGSqD0qemyTS
JlJw8AkuYe52odqKv+7LiTAt0jd1MOORIhY5TgaYVCM7mvgwQ564iMVU6wxp00nG
LjxYmZEBZu5mw1z5azIle74I8LyW8L7kysILtBDy+cnVZ06JfyHmixpz7PVe6aZM
X30OJAHda5RrfdxhhY2j+FdWy2K9mrLuc6qkmVYYAmWo+hwwfNcOrZfrir+BA4ll
ECRCDRYIOrF64J4cWmx+cLdqS8imivQHU7GCZXg1OxCAwgFCegs4ZQaXZfmHgp4w
iuH+wltY0IXvvsO4ONPp+KQHwji6Ad04WtNvEE3vAC9jQ0hWsT8LRpP7Hgl7F13l
sUBXKCXHwVSp6iMGpZdmquVI4X3GtZpyBvku0LF68eIUzaqUcRmk7Cd5RT2HeaPm
9AsNiFBgoPj03g/YzdIK4UvuzlRGXMwknsqAj1Xp3TeV9+qs5yRSOhCRJlW50kdx
XvNeSDRBpDDvEKim0FFd6sQx3JH3EO7dKRfSuvQCHrEAvBo+mZbaUfU8gd6h5u4C
9l9YxBZp6wnPuaCz8yx8DKaLNHjvwOWXh86XAG1p2GY7HrejP3sSo8cCgqcBnl4T
JFGyzWMWG+hVLK7mxq6js+7yHHxt2e6/tYgTuUuUSQKygjw8U/kIV3uNNtl+NtoB
2zLFyvZcL7regchJmYLakXWjNTN76ygPORQdJJUFZSHY1QCEG7Qvbg6cE8POVk9t
1ghy9aZ3jTQATGNUsZSxKsfX8mUYRiPbCAkT1DVQBkGLNySC/vUORJyJEp8I69Tf
Q6+c/nldmFreLcDt+FRe+WHytFVBdkr0C0Dduxqk8zH051owJuAhY4RhWty3Gwok
zCfholyO3IjDCs1zLMfV+REdnzVNK2du19gihC6JOqoG7gTj4Z17GvGvQpqaN6hs
wD/0nPskJv8Z4nXa30ahmUQvEN06JET6XzzrmR/GhL850IFndmDWZqNAD3z5cRhR
ubhqPUp0Q5HWUYm3zg2+urIzNCnfmJwDWs9+BBz0RubHU2jOxhiK4rNg/SfgwLT0
J+tg6PaG4nZZAH7pIMRz4KB9r9j+/vXieywI4Gi+6uQdWMyFoj2exT+j52T8mX6u
iIqOt111rRJJaOjKP/6WQ1Zh+30Ir45pHG+AlsqstL+Fo+LA4YzhIT0uoToWxmUA
i5pXWES5ZisZYeb1gHP15YuFmsFdL9F3hqIx600lL+W5rWz6MIXbMC9DUYX7x/dE
PWpvHcTQeu0xrlMsanTqac/T6LRTZOC0J/OPewQ6j+7L70J7wWwxXH7YY8LKKFVE
WmekfefY0vGXqFI77AX6TW47iDIf5qoPEDm9YbZJ5ga98MKkMHPzt5U4iHxKnphS
hJumYlkYwnIPiX9yPU8AHTVBwreyB+KUPpUuIICYKiFVQ//OZ+yfdcsdJ6dvgE4d
2wu2AgP3ZS8l5AG+lRwJRjKgPgUfwXyn7T8Q3NSNVQMLwNoX7vmX1k8B1JyYjQdo
pdC5x/0yor6j0wmAy7eO0ah5rP0ZaSz9ZEx/90x7AMZ/fDDndYWHZGWMaI7CI0xl
odEKQQILjLgQifkUb0ErchaEILxahLn1lWAXNjNrlUkbe2JsO7pqu1KttanPhfz/
Bof27pSHTFOnOO4qMAaHEMLCHchdyDpK+DsfTq6JuQN+lQF5JLxWRM73Aj9y4aEY
NIRiomyJeUGgo3KEaxKSmYXhNF3MECwlnqNKw3IyOt3Sk4HlO5AYE+vG15NHdCwQ
8lHkMQ6NYEVUefNK5loDq6IF51PXm1Mp900ezHf1DWHW0mQE1j14+E+I1oBriIef
HnHacKcceTHzupTwPF8IRiBN7WyrL8MGFEhKWN7MBQ7gRT59UB2WKPEsteG0bkGz
1RMS2YWRAA8hDm8a0oHwfxruNwG83UkWGvY65ZVVOns3HrvS8iHjP7acCwvUZdR9
jMxPUF7kNP1DOVPScWqsNs2tKYIWdpLrqbsM3f5B5PqOpx+J+cLCXjD3WjYDsNBL
IFCXfthh+58ej/UCH9CN5C705Q7xIt0quQoarb+ljuQi34JFVore67LrCn9c9ytI
7yStAoTdMssR4bzRck9P20dA3XQPZQQOGlA7CJHfM5zqNGo2bU2RWwz8fYkaP46i
uZYEY48F3oymjXAWzcXdhcZ4xTGCiCLponz69gaZ0/5LE8ZXYMbWWwLW8mxVywsY
hVTc4Qns6OkhYmB9J7jJDJhez/uFN5+LiTA1P9U50Wcr85tvJ5Qg2rWLvL0Qhsni
yau9o2H6r9c+2gd9pKmc3xiiLPlPj9agRJIxOIsKc/Wl76o2kWCKw3t8iKKoxlWd
f91q5uuQlOHAnPF7bdmRlM6WZdAU7dZRjLgiAIb/dqbvx26qAi8gq00lezmIH0bC
+GV9jz9lYCWeC0J/Zlpl8LysYIEZxqWV/l6AFcwPr5KnxecHSTowWJKtb6LxJ2zD
efJBee2QfD59lejKwyIXpYLNEeJ3u6u0Ex0tZY+KcEJoa32CdNFVLCTGXzSjnmvm
L5+b3YdzQFSQj4yaXkBb56YhJIBqx3Irdq8b4boL2z65GtIlx0otqXOghSwv9Ohb
d6oKp9S1es7fGP1EEwaArFI5cgHxyZguUAaK7vLWnsZUUOEKpf4zyMsG5D6gvjjN
8sJUWukQJABGRdRoEVuCHJWmg7GDEOv4+aFSN14h88OeR/EnRTdeRpM3HAb8jItx
wLy3LgsmQIWHCwXcTokcTQoA8qg5mp+o8oJMy4qI0OXjZyVz++M3CdbAAw1keTam
NJOnOi09F43qel3ep216AudMogaDOb2Xp1ApNSaDThcG3bIArhVlI4+4IYw1xnnQ
vGc8QZvi8VA5D9KVXF8pwPSuegFpH0/vpUyC9KZbXlT2nD9MVe3oNINqIkSx488x
+63FvOoHJPac075pfzbkf842WCQd6JKCM4i5s2eqwO2KtlFTyPPPB2a4OtV2SEV9
LofsF5qoQKMm1kCsL3StpzRzwWSPcILw8S2Y7KIpKaDLGvMv6R8aNI2lyuCJK/1X
/bMP5mpNI9xI/OHFY+XBHXlzg6S3FH0ynB/U5HKBlzHr2ktLBv1VXALk7X4vD3Hj
ki2cPtWMGulqn64hMnckjjbG/1wiXzV6zH6AP1w1iCfc6K5liaiLsIn0ansU8gj7
Qptb6Mu3XwP1mT9BxtnvKNKHXh32jxabe5XjeAmNHqZebFEBM3Y54T1Xb/w3wXmT
rTJDE3VUdd4ei+S3ZVaEdGb6RsHifUJMGjan3GrP2NzG3Ge/+257pZZaMw5gWa7l
M6XWd3jSahzFaAwmMjtBRT5ZMU/yYpJCRs389LnMBCD6qq32wk8PzDHRyicacjYO
KhTBbUhNJhPKp5tuH9kYg2hVtpKECcfYeUvQ/FkPGGinr3qSaNKGhGsLVBRSVnLR
ex8lexN6w6vemUOhihJC07x3L3TyZohgEfBRRKY7xZEJph1AXt7vbR4jRzhcI97v
frjn7mCBZi4dDOT/GbbD4hJxcTQMvJc40OiP52uPXPGv7xwhqaPxK3i6L86Exv1j
Wt2ljlYKoI+SVYx8RI7Z+4bjgS+poZNcK2LSD4i5y4t0+sojlKt0nwHxvcQwLBT6
najcOAQEzdmftczPEUxIdgW8rMH9tELsBJoqhFSVIO1KFVtig++4UOFY81/maEbW
bOpZQuUatNxmNzhMPsusEBq3Dwt6WFMyBT6KmA6UFseupZKkPf8/BdXM1SlA/dQB
nTorZOkyD926BLDdxtsoUSmPcretYJSrP07boGEJ+94Pw5hh09w6i7W4jyA8W30E
WBtFzG+3+SCOPCf0za800PVmDgcEyyMUTpwrVxyuRHiPbQhIzeoMEh2IpzGWw5Dw
SQtS198aLwPUmSbdxWvVc8xQ4cEgewJf+u1vVZJFNbOhWHn92eZThe7kDJqECzx+
MtkGui+bNbUIht3I0uUPgqNzCCsk/1EebAw3y71B187Cweb0ruovzLOG2kGGZ3ya
eMBVOdzv9VW0Z/m/HZl4V4zH1O6yefdAM4/DxB7FqM4Kt6uTIJQvxO8LqJszdRHh
bb3C0FXVV3mvsntoP76peUCmsr/XXr32zfzsZ2qugAN80lFpRj8/zO0DBTptw/Zw
q1ippCFh3//j9iYCyGTnNcXe9H0+DYr1lRi7CJl2lcUyZt8bIcFriCgz9eiDSEXF
2GcRaUImJmA8JvfY5EdD7BiZwYRdWszic4VEVto/+sBb8ynLyA5Xq26rVhJslduC
SVIUr/6bqucEzAFt13EkcAFmwI8USCz50FqzaVcOX/OkXtlHwAl9Lzmbu3UHTyFT
0jXJv3xTrgdMzxHTBUm8LQEIPV+wbLvzAr+Pni0ZvHXDNNbeFwgEroySD4bfPsRU
sfOaX2PI2Fp6dpAC2qNnqCaexWuK5DfkXu109+1dnEPX2NvKQYzXIWLt5Ia7oVrT
NASYLm52oRhQUra9Tg/GRDNTzj787fK3PUK84M/NquXH1B1Sk7pzGs9pWfi4ueK/
GPakMJ9bmk0mzbhCj+sNundcphqWes1uxExAOWKJNghAkrGB4oD91uqCuIqw5X+i
URS8bXTPXGBYj1ymEqYLKLAmSIzdvszBqicPhBD9veVUlHy3IB09Vy8oBroQS1/c
7xw272GC+TuOxriZ4k2uuYGXC5wZ3tNrZqNtc3nvUzHDZzSZySMrVhn+F7/WVWJ/
xcR8fczWie1kWVpoM7mvCEfAJ1XvWP+MroaVuZCLNl6Gr94PPA8GrW3yHnqcaX0l
VVrhivXnbS2Tp1qMJ/PRMfAHotM6RxA/MZaCulRb1IPoVOgj6jqnubhz/gdpOcLC
wDTJ26Jr9Z5un/10zFmEAKp8dYFYIlp0WoDRrhOXs5tivT6biXcM5vDRXp8PztJX
8FmtI1+nFqcOS8hRC0WLNfTcA7wP4yOjePsBOAGtND6QSRMeDEa3wXBXDnct/lI2
pb/j6/NWiGC3H77fOnf6D/0HmEYvZOrM4fSXQK/lUo0+izieb7OT53sWlTPPQ6YY
fGy8Xs5HjC6iCPwG0bFsZFSdzhou2js7fhAFcJFYAL8vWySPYDDiaEQPxP5HdjVO
LY+yJlL2rEXFvF2Ov2ToDdYIhZEtW1E4p8h3J+m3JI3sohMj1m3KSFIcemyc8/Jp
seigL5huBBdH9uy6ixWtgxZmTRaR2is1l4q7ObADh3qyIqzoXLUmxBRQZO4zCwsI
kni4xNkrqKc53UwP3/bDI7CEXNEXxrjmpMRUkVCSlx1SHzsFLgB4n56WdG4gkRxK
p01jtw1E1tzxLIj/79Uhse7cSrssxnVpnjQoZQ/DiCkzO4lxfeB0DVamORmH37VL
djo4gLczHJZgjB4pMzMpMi3wlCbLpBdVK6oWTdoLCGkVAUWtdNCPV7K1JPvijF2Y
Sabgx3E6T4+CTAd8424XMU3fsL3aIvzWrw4HU0xEuGSNjOpFdMZTWuPkTXeMCVRY
vHKl8AxHrWxOOM7+UO9kFPL6rOjXHdajyLigAdC6KWGqkP0Z3yLG6fh2NuIrKK+P
2RGahwjGVqkwV7hyVMtcfxRf0Y3SeUPUn0j2FfUW2AjKansU5G2RTrls6HXKYDq7
H+lUbxwUz8+Q08LTViY8VztQnQJjKCoqYW/NnSASGm8AiACin1rg37lHu91gyNSY
eL9c6nrQk7H4ZXmWXG4MyAaGyKmaA2eQshc78wC2ekcy/+hOZWJOnu5DPkZ/bZ8I
/veP0zxLImerSzU93Gr0eLNamvszJDNQyVVYyTcqOtJIercFoMIgIp3ebQAigkpx
C5TbcnIDbSHCYFXhX5RGtrHdPo8t8vGKcTKQhsQiqV0Mb0xoua7WX2e3H91MJAqF
g3WPK2t7AHshMDv7q0Zi/JIS8RuEk0Xom24WkLb6fIDO0myLk52E/aDl/D9ggOFo
ocrF2AogGpqSI2NY5XulPFeodphx0dz0ifYZrx6a4uKG8yHcWpzA1VHUdl1BDcMv
9r3g+ab6Sm0/c5NB1zq572o16SkTzGZAMpDcFOooC24fk765+qAZoedj6v2gxZuc
aQoTZcbBke+l7YP5NazDUAiOILv6pBMzmnLDmErOWZ+76zn90scYtyiDWVN41Ilg
27DqaDSbRkpldKabIZ3sUdqO4j8xqio6ahz0KpMJyTtOBb1TRzoG9hrNNZuhPPpG
P7+O2Io39wUL5E2a6dnr09xwZRcMjacrI+UW5gaNtZcwgclLF9hxCJ1FcfrPge+L
hxtB9VrAvsk4U3FXad4atP5cbMPsiSPNrkrVShSo7aU5Iy2JnpJQKWQ83Ero2LXx
BAjC/148QInWOwX3GIkMBgqFy8K21GqtQu6Q162SdkJiZ9xNiITK5KqRQ7TIlsu/
iXhD+HD3bLs5xGuwWi4UbWGIIdyebszPEt7zEJmJyARhYIgjjFsGgBJ5zbYjyG8Y
j1xTNDa3iDl06ThY/vUTXJz+4hAqD/IloFS4U4Zlf+/4/Hyxw9XKJ2YtifX87nZq
M4uwdm907eFl6S3YGks1ohbdm9ts1GN8W0A4Vw91BWEFzjG2EZSm3qbC4QydiYI/
336xo4iPPcn6ubgFuUWRv9+iF7/y8o/UEFXkAjZxzMrn9QnGLzbHYFOiya5MF5so
KgCoh4FoGn03LA3NSgaMzhdiZGp1Vh5sGcuKwtfQ7Z+U9LjY1c24qKzqmzIpft/x
whmLZNolS9qnJhvqdrc2r0D30fwMUIZfq8kR7E5ccjFegyuxrhfESciMBPeTl3u0
z3V15RVXAANMF8jZuKC8kR6/9kUXjzGeHg1g5KX6O518s7Td3Inuoa3DWPpujk9Q
7RNlBSAu7eqzuZoxJtAKZ77vLhczjtWM3SQmkWvTANWmAlSMrpQsb+FAx5qFr97/
FW2w39dsZ/sb4y/Dfz/ciaN3Yr4iFu63e2s2c9ogAZhVyO+fxcb6kjmHOeKlgt/1
yR8Ffp9BqBGFhqqUHEYBizhTXwGySN/NeeSIX5dJM6WER8mwp6yvqBtDz9kZo2fh
FIFPmMtIVOZTonticjTh8TUzJhY0bFGmD+/uA2+ikrMKu2c+zHst9JVb/CBeIx7X
rIveEPlMrQuhzfg7woyCM0YVc1Y8TCB7E8bY0qru0+wWwAiVQCbvseqhDTz205Um
kSA0dRSopV9JJsmdB3FKYW/4myDuZQ5HwljXP4d0bnHLl+2iTO8MMS0FJryD70BA
ZsZOyRbxAJtJb8CMqCUGeTi5bCMRa4RZnZIM44pkRsaH1k7Gor48FZ+inV+k1E0s
LyHepkb8iQdAq9ErRsKlhEWvU8gW683CVlvtjEwHa4aC/qbr6BdsC08OASjnCy4b
8ECj0uHYZHhlYvrp8EnpBWn4RnFx9GflaHWMVZtt2jFRBQ769YGp6heoXrw/CsoU
k8+rERQBbYxNzGW5j+zYEX27xqRkPmFVUGMbT9xEY+8APVKHD85Ntnlz1p15wQio
RwFmzl1j/YjqibEP965xCF3qKmSL+1DOYMbblFCS2JIbHZc/CVw33jHiagdVnoTn
pJJwyjzM9+n+Kx56iVjh10deHfiLvyy4JxiHMPY0M122UaYuHbgoqekz0JjmviqZ
DXTpgSwtnkvNLBkWsbsBfY6FLIYJmSo9q4y7iC50+UEMm/cgovP0m5TnK9m4nnIW
kx36RN4lSPEdDSmjhF4O3MX7HMGHpugIanfdzVvP6/aKA0tiXznGus1mAeBZWUjE
TDVmo1du5Dso8AZbR1fviO7J0+1x4d18GFsSJgnyT+vbJhqQNNTuaLAF1C4wLpx0
3y9WRc1Xu/m6vVUQ5svuGYK8kSKDyV4zEfr/VgtE1GedIssDnUZfaZch/fWM32fV
Wdsi91VmvlzlIteeMpOzPFWR8k8O36CHMxvrRQ01Mi4eKDvVGqlzJeB7pVtWNkiJ
Jdudmzeb7OB+uX+QFgt3nZdjOJ18kN1iwQhtedJphcv3CRa8GwN7BY57RZvfHTTi
/sOGXWISqYWVmIpGlp54UqQ1orm1vNqaqQ5BE6jtOAVW7L2RbSqRRCOEBPomMMTw
kLBGeYGEgT0Jy9oyLjmLSbwaMH70qTeYN5LANNLNfFKom+zubBFFpGuhqltwsEEU
MdeduxhpVdDl9Oc/K8KpxfPEl3hNoCc/FBMOuqwLKBFMXXyXz49YaZraxZrFSMfc
ZKTRH4CSxUbqmwRVB1ragIWIS3vIJxF17OoptiQKzPX8LQe31ngiC79Zkk2dAScb
SvZKtBUO+5yYIFBd3KoqWZkHFLKz7WpNdamzIs9RxdXyUZ/Wo4E4HorV5DMPcPGn
JdIKWD50KZlgiEibIKnzykn+jLj1ns5GW0UPppkT6vuEY0+njppYgj4VadKTOKzH
CsTPp1nW6FNtB4Kyf5DwnZIFLcyTMOS3a/5P0VuNW0vZbCzf/Rbfw6yW3MmrBHUJ
fLHDyGDBGSzYS0TOluhfoQU4FyQWHiUTpKo4rJjdypTYh7YA/glOIlN4fIBTsrHC
t8AfLlhOslhnhzpYazkqx48cny55NpWT025roPQoAyW3NoUxmD6g3qz1H9ChuupF
nUmohD0WdRd0ySp/LmTwhufvP0/pMTjCayuCKAMkj6MpsgNXzf7OLIFZ6KmjR9be
rcNog6rIGvYqh6V0iC3Z3MxspCxdApOU/5nTKloX5KvXvgKt4oSipyHnoNXZo18/
1jWZZ7WRNEZl3PJX5qeFwcHvHwUj29w0s0wLyuFto2AtGm7tR+ZQxEZ/65ZO7bQF
FSLUiQOrV4S8uhdKG2uULeaIlsbh4bTLtwp8hFs8cYs8MbTRl1zgOiotcanTooh/
zRjbmRg1TfOzM+9OeiU7NmZgp5HEXreZD1x2DOh49KNdhQYmTFoUEAR/pBSnisD5
ENTWnyN5wrj5LdMCP7nf66gV5hcKiO4DT30oQYoxYiq7FMK4z6qNaRAbimO7yGG/
JHnB4/zFkhVGAW5wN+4ZxXnHrWWrKAz+Sve7scB7WeIGcA4kxoTnEbaAV4B8SO09
ecc6f+GWsOivFPyypVVSIx7khZuAqUSC6utLam+m+uGaIR3dIryqzNHEQABTXq+S
2jM55ZYJQ9v/NVPBQ5r8Cl1XR8XRrkERpDfc/NX+bokb+Ox6XViMtGfUBXlaAnEr
0UyjtNbmQHcWiX9bKp1h0U7Py+j93zgzesd8F5EKxufXD79wUEHp16Ec11+NxJmD
vMl4VJyeGBYNRV7DLY57DQLlj8TtKCm9O9CgPN/rAcD4CVXbwsU5470bCDI0QIRQ
YwLNq9rTQeaz+U3P0X1m0j2D78J4Ti+QJdiuj+IpV3ShdZ25Zb01C/eRs+uxj9rj
VbMBUu2vBhyeMG96UmqtJniNYrs6iz3W+uxXTcUiwr3GqW5jVGFqmF4BgEOsdHyB
65CYU3RvaqhwFl2NDaZw9NVqUCQIFqoIobRXeh9zOr5P0HHVRr7AqL+iDx7TsjK7
655S/MK5VXFzW2AKvr2Nkt/qpp7vuQn/jTVPAjVqhhiQZAtkjambqiF9Q0VJDVya
B/U4PPVDf7jXAFW/D0Q8atSK7QDAThLIo//ai814m1Wj6rNeS6Oiqbz/scdiHlvj
58vexh9i4JGYp9ZcfCZTEH84xymAdoQKI/fNQ0rJSeifLlun5pqbUD0t6quVMzO9
SvvEY/+w35sK6vVXrg1wzgkpIc1BlM4JnvbW0UbBDzZghWomU1ZPi5Zla9y9Dz8Y
8mxjYF1XziOhr1KQPaE+BRJUrDWC/RZ24TTrdt7eF4eu/FGkyqFH3SxiAGQdlQw6
4Ar8elZ6rpufHiOKkaGJ1+h53cd7f3KdysLdzljldW4iJrgHB9Piq+MbkbHDjhsy
hNSkqdtB5LXQTh/PdawjFDXP+rnfFoJ32xQDvvqUvtvziwmwk3PLeOYEQt160qmb
NlmQMFCHJ3Zajo6G9WnxqwegdpVfzKTuYpVd8Vw8sYu1HYDVUrr7ukzNZaCKA1D/
P0ldablUf0C+thzTbszLBxCuqxV24awum82UZJXkFJyFV//Nkz7q5pmSpQGy1eyC
5+3YWupolB2ZUY6DJMM2/aKRU47iyId0Q4zqUlOI5xBcQUUWFoKNLZZNPHKMK2HN
77FR/1J17+t/inoNGePZkb+WkA4DTt4FtLRP6fQV8ytlNrkaK0KLd3BOPuMkjcsI
yIzw4zPbepUEiNSePVmN7cY/zytoiW/1BglSxcjTGMXO1eIYEcB2J4CtG7YhKZu4
jFy5iLZe3HKSbW1kOXPwR1t2HvIWTD2GuICF45Ji6jDe8RyPPBXzv2b0rInYjk/1
Cwdl/8FJHqwNb+5P4+vhE5D0PAoYrdMY9l85uwErwfDhT8bA1hLcJggUcW2xrIx/
BjCiFy+ngfaItOYmuRvTiHt4p7nZ4nNa1qZNSjsh9Y5nqXecHEuv0rlg9qyW/GLz
CH6P8BYcOLh1b4HkEsHOTlpAzoS8ZHW9ZmSIig0awOTrdPcbT9BQeFxyLtL/lX6j
QODoO0+3nGn7AmTYy38EiW8b/uU5RBcpHiJ7qMBu4BOPNL7XoMc5Z7GYXjOlnnIR
SOw/oTQKUq/Svrpv3ZcuS5C760JSjaN1jNydp6tgQsaUtTdtk6PSRq80+DvRee65
qkAYS//C4biTi9KsM2z6Xy/SZSi/zchCcWdiuGi7j65pWbjFKOwdA6NzGvCt9D3t
MBY/p4wne64LjgZAUyxMcj0HSPKe7HfP9CTIl/q3QHLZPjLCeMpUtfiCUAYL692n
sLz6LZCsOHDzYILT/oVs69DqJGCE8RtmQ1TLfPkCq3R+e5dOmIZ4WB0FfZ4ZsqDs
cFKdmRa6LLN2cabMv/xCHGOoiS8f5zMCV1nCIY0X1Mfp+ihutY1FY30b+e+jNA2i
btFu2z3j9zCiKdjk4G8FRnd7eqb1+LdCKYE4P2YhjRzXzZr/wcGAtai0eWlfaA7J
NgNaU+uue31ufGYGWvF7NfKmnmupGNT7wLnBzooW/id4m6nMb2SASD0Gm+8vHQyx
da23jwNWJ6MkgzK+jRNi9MBm+8KSlLFtCcbHNVt74oxd4UW52PVWdaspMGGdm9pn
FFVRBEBnFgfFR9jBa/EpOhyhSirVeK3Uwe0bMxsKVDVHeG24ItDEpyVMgh8PTCrq
gQAVAwfNQ83eOHux5cUKD8l37oMSVHYxTAOX1domjXvABoPksVltGppfJ0qe1f6A
uHFI3FPjXRx1YAJ+0SLAbWdafI4NZlJP+5S1pEb6inJ9Y5KUtOOA2FmJb7T7DfLO
AHmVI30jb8dcFDGSCwVqX1cV5+lw3nLM+zHjXqPobno2pgPnjXHAHjLqMp+V2hBM
6ID0LdhHwZsTW2Mwtc8+3m6+N1/0LMVIHY6x+i4rygJ7THm7IJa03MZb5RrguWut
gz5rtSadj7CjdJAvWAb1254pax/0Rx/Zzu6aHyB1/JUIS0rC5HHkpX/YZ0pDig7H
ewznSIfxonUdBiqAHjm9traSta1bW33zsLj1K8vXN8FUO7w0wtFRdc2jHvfeiphn
MhereQjj1HvrDz8Z2ynkHQMk68ALI5LZ70FmnznTqdkQNbq8K4FcR41uipUHBcL5
KYP2BjNZ377qtDkwlMbl4tXZThw9eaflldZqe+xbsp2RuqavcYv4FlhkqHggMdqs
VL+ZvS/6Xm9j4bEePjnkZ4Y3Kej2cw/fMOrAk5bGIZOW5sqGs7CYovzP86P7d+uj
xn6q6GzioP3HoW7wYo4FNbHDqPgOa59TFgYLqTv3n9DSOxXYFIDacHbV1L1sFLpe
8cAu45bQNsWB7TUBdwsWESSzmhLpPLVAGtpKmMJ6ZGHhXzokL3dtP5Sppv/dks/s
hBaS5gSsdvP3UP1ZpYcvzbAMhB65CmaJQ8nLIwnZRXqWBdFRRGlO/vnAIE102aT8
H2Ud3eOYkUQyxDAR0mZzTc8vFqA1m/+QILGVuskuC0wXI3hVm/LuITByo6LKRXBe
V0VQeESrLEdG7fjYxBtxoTCxuLjBMu4MmE/1REXFcSHxJDZGmhmMu9bjkhCHcxp9
/77CR+DK8QGky4SVGAlz1zfCFS5EdAR5p7kGfNTA5Os4NHdNF4jSQYeggJnxWzC6
TOxCHjjThnlZCx0Aco0tM6gOdiv64Gpe5plVjZYurycxwKB0YlJddccsxEMz6N8u
HwlcIU/OUQQOb8NyMFALH0DTQiUVq1QfCrywKmx5XZkFrA/JIg04w643HOtVhAp8
IWE8GrDVpeph8108Duv2W/og2HD+CP7Ym+MnvGz54mqpoaOEwqZUGGbS/+WMT5DG
zbJeTMNVd3rmdlSP9btnssXVls9Mhtp1K3YGgh0xJFfGMuQsMjg6sNHvxiDuEpVW
JIxVIcAExOcoIV8dLcpHQVeIJ1XbESdJuoC800uYfgauTRY4nbS6fx9/pVsqkT/F
WbCrLw/a6R7F+8Sc0qZ34PYnPMRZo6GM43M0bM7SoiOtvkkTWdlTRTCCNR4sVE2G
VVCgyq0vO3b07ldMNFbEYNC2ssT2+jzz7X4HyOv+toasNKBUrdnqO7aSuFnScU8B
KKwT4z5gw6A62wiMsxoNH4Li/Z1iJWLDql9SfT0Tc+/ElE2J6dsMfZ1hP0pbQOR+
ns4iTQ9QoyCVSzGK+kOtCMufhCA12tteo0f4LrW7p1HjZ+tAE2Xxxx/9/mB8lmfj
8DtM1lg/Mx8fwgFtBetJeyJczn7AtEYVj29kxv/BBmKuukzKPY5dMSoL1inJSRUK
kBou6dShg2wHBY6pQcrBe5pNgDH6+BBrwxsqv6GTQP9wq9NWa00UfSAMBT2nKy3F
wk79/V6Vn3qW8qytreGpD0OToFI7DIg/VNVKHN47F3E+S1AW41DrwtWGnXJEyPOR
fxutRKqwqPxPcI1mOYDZQlUeCtpawT8aYTzQaN8bHi+EO7H9hhEjiVUnUssOSr4i
UUeFtGCYXgiZ+2s4ypOOCtV5kMg2wJHm/7KoFovZDP0hUQIC6QqpmuKR8lFQzfG3
Y/B04TlO5Ixc6X7bomHzDf/f92OkVwXd/0a86oGNnlv0kmiwPQVnuw3/D6aLKe7L
tOHMKtI5t7sKMc+aOBP0pDJMqqsbXxyr3Vwk986f7WG2gllwfN/edqeN7rDQplkN
V48Qv2eVkURAp4+6uY2J4kUob6bKRjcuvqKrrILAAWFehVDJopkAhQ7o+YRQ0q/j
IOKIjPyRS4nEXFwifRFTPm4t0ezWeLh5Yzw0jaNloY2lB+fW/RvgPXuzuaGqjXS3
pkR+weClAml/uqaTVDcuyYh2SeJ8gLeS5XopPTlox2abt5gn/oAm3lFAU3uG9BGd
MDONQFu9Nkr2FFaqY7EuBuAsuCClDRytxc91ZPF5dmwUPFcAnfehmRG1VEXb7zbS
MYKrnngU2Izbi05+RzblOSwDU3n54j3UBLH0nWAj36HZnXL9k4OVXkD5W/Cb5j/J
mf/fO4/Ir8VNgS3GjZMaB+9Pf87z/IiHsmr/t0HW8K3u1baXGFM2YUKRECzCN9vX
uViUI4eWIoi4lRxA5lfC+RkL3o6LlmfFw3PNWuYKbVXSrvk1RDQxSg0ViYQW8GKr
lKaZ+SDOemQirZ2aQiQ7Wg9KLfOZQjmMTiFxP76VbrPd5bXTBb4kAfFHP/KG5xs9
bLS89stZYsTBXNDCabjXeyreXuo2Sspx3vtHotqu/bC+Jc8f88Ypt9qDNt4HsjcY
yhzYG8jKNZ72QlTaCp6b3+wzIK2j05VdtqYejxJNNtUpJk6H5d8YxGrhVXjNwpf5
mU3oN2oYpdVQTiC6jQyoksxtkJEY6VQn/cDSwW4/vKlxYuDfdmnyU2uohRdQ9o9w
E/M7HRZ2gz/PvlMW/1Dj+GyJT+tyza9pIggknv/Y/IZeYSAtU4G2qwijp4dX/GuB
Q3wqNe40NtUmpjhLe6mwDBxZf3iSyTsWTdXKW+YNks3SOv2NRA/QIWTwiW/EPW46
/uyDy79DGtmnuPcW5pkKxNusJZrMgt4f5xCI9PpwsUpDhNQOU7eM6y18FuluK2q0
zMlnz9WJIj3spvhliMDL7VwDXVODIoR/c3UlkqPLHikDg9Lf0J+FvmQvuoV3DZ8s
/i5U9bz90lfUPPHylyqtEQA1kdX/zltdwjfl1oDdVs8QB0Ct7kHzkO3yA/ZalkRO
dNwfgUPAYva1D4sf3iX8UkQGOLecu8aLlQxvkYr/BNvzvPxJw605MVUyyLdzb65X
elE14BvFUufu1zrZjZI0m3b+Za3Gz/7gQ31Fg7X1SCcvvEk153SSz1Z82uUsEeqv
9ZfoxZFS4LdFQJ3ZibZ+x+u27vFPOiR9I9INidaVB4KdurY+zd2dFyW3Ty0mgt2a
/j4L88gckbVXBmzVxEP/irZygMzIr60iVzMUvDVkV4PZDIkQMg+pi4iB0T3rt4Q7
6eN/vdTCS93pAqWnPrEvwEvbYuroNLE8nam6djGd+myGs8nOSzFWanV4O780AaZ8
2ewf6B3s4KKYSaTTUItL0GJlKzyHfhASfhWJZC+qWd/1uqHVPoy6WZ44me/yeV2b
Fq4S17TLC2lPYrU1WxNAeuq5goJfwN51VRPvzLdOKSosTYDXHLbx9OPJfWaPpDu+
zDDMXT06WbzEDcqzhsxh9DaUHGyWBFNNAUcVizpskFEo1yDqwUEg+CPc/DuZdzRm
XxQqM2GWp0VZTN+2jBAx8oSNAGbdB991yWT0QK0YDXqpPIkYp1Hxrk+13YWsJAiT
6DKtvsmeBMmLfu/fs4v874SG0qugg4NNsCRmdgv/jmOBnfPHprxk2FKBaYqn7My4
+br9tU2YGJWuFaMGJVdUIFLqfwyOS9xO8jZXjp5aUfmBnU2Ca30YRoLuhO404J8S
A+wWYoEZUEI0ROVaWlVGsuIefyenOnFebYPB1v0mtldNDzs2+gE9OPUIz9U8oAP3
D+SR/zh+qgXhLFD742AKHC2GvqfYOT/34Vwi1u61z+I2xfffxeQ7Rtje+kl7f490
rV95/EdRfVw8gqeZVMtdnqkFDsFRmgKRq1mgj8T44Xt3W3lH0css833xCCGOrjph
+/nSN+t5qpzP3QNs4hGNXRIGG0cKfs/caQl6mxOwjEri0d8CRhdHVvl1M3/SX74i
6hhBYJgrHQRsm8aGnz9X4T6q3F+keufsQDcnUzujxsYcfI0xOMDw1eBEJ0rEwtCR
mQyeMFtvLEwyAyH1np56MF9FhhIp9c6oEpMm5JEDclWguWy4Ek0XQHj2Vrb914q2
Cqhiryxgh9XQAX0nZkRvu3vaYj9TzmYCYFa88VXWfIJwUmz/wVkb3C1u7iFuq3H+
hSMWtBQqnzXOIRbTODeht6S5Q7Gb4DzTqA7r6M2m6W9uYsSp8uanWt7Op4SDVaIu
2EFUm9Y2oAvq8FD4eWNMEz/5MQQOUvBBjiOQanIyMK/HUTAaOTbgyqd/XQ+Oooln
hSHWKHpQn5sahdBUfYhL6ajK/4Klgytz8otxGpHjsp4cidCjdC9wn6UpEAva1hzz
tFfUqRuatNaJHi2WGKdmlHuy3dnTZO7/ddUpfXDZvifFGoer3psZLmnXLdHmzFvO
dsNQ8Au+1VA3dBrpPzF48hdN2rgfRjlj7b07gAIG7HP8R++NiXFHDaPG8H9sHqbT
UcO0ZS7uGk56FD24MRb0+Fk8OzDXsKNTYow2MSpa9Lh4ieXnh6IRuSJcd6FUJ3Bx
nFTcmFxd8xYwWt0Z8cVD6gVlyS7l/OFlkykpyBubcoxiawT/8X04Y2LLa5Cwen1i
8mNRWhe1Qrvk9AQ120YSrvSV3p4azbh40Mpa9TDDWDauoyqcj2g/ewDk0tHN3DHF
xdptB6a3s6UhmRNaIgUiJdB+Tb5fiAwG4orHGS/DCgzspqEUl6k8Zri4fMsZ59Re
F4a1EOpRRj4thMxJ9k6UcpwQpB04bOQmH4s/73ZpA0ICFPUXF5CKu14HDjt0eYyD
vALvB7awmGuZuoKilyfVrZi4Pxho5WzUeWW7PSN5vuCNVfUD4On4d5eIS3kjOA6N
0a9bS5EwD8Cnvq45boUJ3kqMpNInugsEfI9xJC5ZDUtDAa1J/4SZOAn58ZcPIWt7
/LDGzjaPK/HdI6rvLgLgr1+XpTeNNWl5/g7L0plqjz7CfLtxVs6/PZwsjlMUKrga
HlTvRCF9FCp2Vj3rkimsxylhpM1dXFPoiqBMrsYP4de49+fj0gbqDkoOkumA1XR+
pZPm0jaAYfnx2WVvS5usf1uuFTahS+xz6VkSpGYTsMzoo1DQrV/LKiklfaBYWNp8
7GGUcKY5kmfPyvyGwaSUlsQtWNQf8rpn5uVr+TtHa0vFN1ebXbl67Eb9yhCmZPJP
USQ+E5vJOz3J2nsfeY4oWWOPLXAeUIC/DEtAORWDA1KD/rJTYqw6PF621mnuRcAi
B46BtHFOqx2B99BPXJys8ki5AT1VB6IGE/k13+xVa+NAvxF52HOgo4+UqpThyfvn
wdhfwE6DAW9Ta5cr35jbc+Xe7Lu0iM0M9thXfmX8a4zgyb1AYwVsthbTSvmvNNm4
mE4vC743VbGDJfgmIGabRMEKldHSQK96fYs9mKVuTZGnGXHMrxrCOKJYiggkBgX4
m7n3vBdj7+exzxzn7yCAm80YOLaZy0OKjEahmQCYh5N226m0s3g7Qts8h5FyxDDO
yWnrIBv09ihvn4wgHQedToaTBBoqf1CLtnZ2k92e2MIj7xt4mGgNs6MyUzNwyNFW
RgYQ5EjEpQO15dUj859Av860acG6M71vL5XEVuKphPsr1MfgcvFsTwddp09+a6tS
73H6rwgbT9ycgybAXaQ+HxdaWsVLJ+fT6f5VJK5TpKdxOC5eGuHfHBI+Qmpb/J8m
DBFPMYR4EpViUGoQs2C8DBaYRM/UywF06nm1UtvGfvXDmKYu0g6BMz5rqjJhNjNd
L7kMKCurgHOQNd4OYj2zUR5KBqbFZ++lT+4xelFUGKwzU5Oh9D3r6sKmH0SxTp1q
PjZHLgKi03FDAPhT4PxdS42SrKvWP68/f+sKhvqm1A9Rb47y3BWzY32GnZFMKFWR
a8Ac+aMqWgJPHdcjk1kTVHd8UbrHZi6Rfw8YbvATQcZFn3byAKPST3rKBYABRemp
1HLWNDgXyDbmsV/F33RF7YNMlCjJ7R7jHtHIhdWLjUgl46w6RG1Jv6/qmlJP7s3f
Fb22A/dYyUy+d8JfpQa6txmvnBzagY4kvIlemc902MsBY+PObx5PQhyNamCpGAex
kkiOHkodM6FxlD6MGiVg6b2Df7lTSLob2j82d6VWhKPFQ7FLV3cVqubMl6/NP/VY
PaWFmueCL6IlmIZCe/RtfTwBQvY1+9CjJhRAPcUWvE6oUIgrQIh3MjN4fHrNqYEl
Y8ifDg5hqUGLJag3kc2npabfhw1cQAe5IQ9CbnhV1kQEVjX5MH2bcFoXlwpcB5N1
RrsGXkozg3PgjF37oTz90iSmNGfkr3gvxBGopj2RFvkJaDGSHP/slVeEOg61q8x0
JOm76TAk0FuwtXUp5v48w1uDgFtrNPa9oq+9smikCgHUzB++jeVUleyuU1pPWmG8
yaQH+xXjnhky8tAgIZ6zPJx88XP0Ijd+3V6Ze5LMDIEcIxaDeGk51MVUTYCMptcv
ggegVSYM2+OpD0oI5H4V3LlLVenzRnFVhcbi4sekwAUOXbKFNudnPJ8Y5rf/fAn1
nyMxJYjgEwR5WrlrqGJCa2eWt6CsgnQ79oITGOs0XE7jksbt9qda1UwDTe2Jxv05
O2ihrUQabgbDTjIG5iWJOT/l9MLtUjmXZHWUi9uQNLoKNFE+1WQNw+H8S83jzKVH
Ix4lYAOmTJHVaBS+k9f26xmJdJik5rv9/nJOGKvjzGc2G5QeMDlI/dhNRBJYBcN1
k77WiuFnwsGwGNEMYlQBYEBArWor815LNs8Ksn76/zs8hIshd4I8oqHEJgLYoYiC
9/S1F6HB0luOlGzRixO25rgZiVX8TcebfxFUupmCMSOQdcbUP3WyP10SvDU3oJQi
rJP7m88ac2z8zhgDGWRuIOSYbCZp1ttI5FrmNx9pZlS/XBf9Po3WQjZyf9ysyInA
3tcbpxkblE9ZPJjpYE3/g234MsGlyNz09BDYX5oZhKUXw6dAZivIFfFen+03diyV
bHACajQwyP8xzsmaQToVCcTezZl20Tv+uj+iNyCZY9U2t265dx5cpS70cp+3Wlob
/ML4OODOI14TdLA2CcPHkuqOV8SQmNJfVgBzLUKUH8qE3eRYXCtJAz3lpgDUtwAU
ypEJzKMxwdqswBDKzIYM/NaQZijQykAKPpGRk4W3zF+U2y9MxniY0rI+aoH/VHvr
E8DFbfaMaJ03jVK3Zj84fuZ8nYnKiUdk5nV12+NkIY3Y6Eu5UepbvDO/sTHMVq1J
NKVEU2K6g+1mU4M6LTxRTGmpSio7I2XGSFgXmumhG0eYZG4HOdwBRUulC0fneQUu
Uv6q3vW6k20rYBnm36E6hFX97K1unOla43yF57dPt09227qAwZVON/SyEJEV/oot
6nPpo7cspMbqXvzDIYIEW6eL7Vn6Kby1QZYrNxBgRHjNY21N5udi/PuKZ6VyuVmr
eI9X8ERKR1SSMg9WHdWdXFCqvqUSMnqGv/C/QH3U3KSJXFp/zaOKGxFOVS+me/UU
1PBqIEXXCFfgETLLzcw2fse2/03VUY2IGNTFe4gJXUD8wpQGNzOuTrM+jO+dCst5
JNY3ERZqFxx0IK6h/btfB+6CqiVlhH3n6sMn6kPklorMrJEjDw2TfOLtl5sWPDS3
PvE7iUUQv1vipJnw3/hA+cvNlUQ62gR03zgvcXtWtjGAhSxmxA7FYrUa2QAg6l+1
v20x/tKe+koKvzek7woUWvIxNeggIUvfFwthekPRHIHSOBDOWsVGFwhg0mHf7kF4
VflriVPk/SNhsl2yWjYSXkDeh0XK5mja6xlVnz3++RmYcsZxpNQALJOeGj1x4Q+C
mLbI7g0IVXnJt26m5n5uucmlkacENs+Lj45kkT0eh9ouik/Tg0OY3ULChZ5IXUuf
uqT3T2FS79ibY3dou8cXer4kUu87pZKqs67UgmQdS+vFxfSb8lB130z+o8OTtiAi
9l8wO6NwVTmdfgp+x7LXGt1btMUy9bEZkl0h5RS5UFkEqzh9KaPO7+dgYrYYfQdg
HweVbiaEUJz83OFALMkIpAP0Nr/daMaqaysqxyCtHZT+rq3vCP3fUPlIGXlpBKZM
yTO77NQE2t3zt8eL+5tdO9ANj4hHlmnCQ/uCYrzeE/8TkZWMuYD4p8kokL+HSl0y
r2YCtAlYnqJG39iNsNNwYBkzRmUaXEsFXunayo2Od0MVep1JeJnI8AL8A6pSSdYJ
9xq+LUYUDtnH8CMHL88jJCIoRy0lYC20eUwOWCoQz510Ko2yfmZoHhkDt8j/gJTU
/Xvbmt7fMw9hX7n19YLZgZ3XPUpLnlYDLx9ouThpGHqa+UgNg3avE6BuOz+S5cVO
j5EFNVEaDtu3PWG6Z/xo5X4W6NFX8L7m3YLjnUQrWJ9avL3l7z+pd/f/1GeYDwqL
JdE3sXOFbHVP8UvD2Uqs0zvATj24joE8EHUffBgfXufEcAjr1zU+TVBalK7kpJ29
HJv6J0PaJqoiT+Hfk3lTSy3LqilwPK3OdtmcjVS3NLdcbUzr2Hsi0Vz6AMorrCIW
VBwuG+xBpuvx2f+AzcunrMSNm0l9+LRXM/oCSf3Woe9GROAw+oa56F7EzH6PZ9hI
kF5CS/sOKCXxJc9L7hmXxKLCtzdo5gnWe2aYRemydki85OjNtnIDBog96aMYtxdk
hAf4Cdo9sxQvrxHSRv/l6bEYGwmIHmFZfY9vQ050YEnSLlRdud3yEtnq6o4SrIOh
rGb5/94jxrYMzUtkLt+f9B9nkycZFPUibWaAgM6dtupbeDzH5kNtsOQU18bm3iMg
ZOQoLU1yyAy9J6sLm56bedu8zCwuk2KJQErNrOrM7ywjea9b6OiqAJIFvSD2HZoo
aQ/CYGpRooY+L+S8aFnmyMXhXMlP1EePxQ86wwfBtVkWSApD4TynXM3M16vmdRcS
wLAd6RgRo8ggslCW9iozBx4oxl9/1aByQhu5jBxGpEkQh55iuEITjhln/CvILMwA
OGhQsDL9dtsisuUHG4sRTy7LN5x8R5A4+/LwwgostkuehcZYJBfN+hsEkUcG5hyB
xT1QilkudQbxiLBpGOtZFNv7jhS2Ij5eNa4Q8NKsiQ4cLPuWC7V+KOIoxzLo4WW5
95jKPJWZn9Sp7UamYT6rXaWmf+U+4s42uJf0p9LQfrvPFo5bTTk6gmL4PfEMqCb+
yGQ2NZAdyIl926Wp20IKESCrPeH8uwMVQGiSTgGqtewfjikroVB9TLyF2MI8nFhl
0rnNY0rIBLA3+2W+oIeRvIgB6KnoGXSrtodnOGaWmmLLJRzOuWeSZPrg6viLVy5e
jAc8pgi+HG/Gp4XjVFCUMr4IWDCgdQA3GAE+p2qRsgsXant7c9VnKuIdKdxneDwu
vJMhBjxpxo4lb5z5CjQKwkR6DHWLq+V9ai5VGMsgRpSXVdFMGSB4dbWimL4aYNyS
YsqNcxaqpe+FkPCMVHCHvfx17VrUsf19k9U2YTaD4iszhKkdaXHfpU7vFwMIqH2z
wUeFU+6PWnYrJCTyVSyn74L3nWG1JsYqcRerTGy2KIU7hE33h738xnHCZtCjYadn
tc6lVxjaDbs3uBUB868ClShsuNQSFIC4wyybOaOFbK3venUWr4epAo2XUGcbdHWg
1s9X17Fnk3WXrCBqON+mPmMIDGovhq99elBvYR0T0DL7QNnjOwtLTu9dmnRvpS9O
4U6AMuSBqFasFmK0s61myU/FQUqTSR4IdL0weAs6YwhuFWQLi762Vy01Ep5bqact
dr2mglz1lHlSvVp/yeZE8pWQ/s9gaW47Mg5aOX5/uprN0HwqXgyIxDXcdVj1/K7R
57tfK2xaJ4AowYpbjqU5P+sTt+eRKSBb4VTsHsNpaHwmt7/5k2LtKuHE1Ha5zdUs
B89pYiXVEOuLEQcR/2eEAoXhLk4vtiHuuqOHCmZ4P2FHV+4AJt7cQ+IEQBJiO9Z1
wJp4cYBnR+XafDzr1eBooGJcuFomzZVCNuvxGAzp+K7Xf7f/zn71QvLKE7OqFBHN
euVUurYXUtHfyzFmyGfMBeCiR5WqFAJLycjGuqVK4ji3PYpgIbty6s2eBThjwjz7
EkqMNEGgEzwn0u7xTyODWQR98j7cy3A9uBkw04xd+aVNg5DBgOlC5yYr3Vhyksh2
xf8IInnWsAZK17FMvBGzbiMowk620C3VRYoxYYS3MZY7I8+uhwrrCknbVTzznHag
9K/rpG9VleLJ9dp4YJGJy3nNdIApgSwMfbSp42eSqJOAagTr7oLU/v4iVl9UL8io
Doay9EhmiQNe6TpeXxXpQfSiQh7wKXD4sIe8f6Ew7RdrwJ6Eq+VbcpPOSQ16QwDs
fjUDhS5rTxGhp148V6PD/h+sDrHRS3VUDSIzrB2sy+OjGjdsj79MlFIC68ggxLYA
2ZyIR5YLKZ98OSB2p4zgJiczI/SodjML/NbwfnvaacgyVApSHVQoPdz3x5vcM4Yi
xkaCe4eEI+uA+kGi5lOXZl1thHC9/c5Xmy7hFHfJpoyacSiIkd8eLIesrt5EM1TR
Hz/xk7ISFJRyqdhRCkcpwE1NIhpdkwObSwa9VTRoIA/DLDPOxXeJ27AdtTWL/hu5
8KP0f692thp56N5UGkrx+sif8+al8Ze2lQbzpHLtCne6YCBfeeAfa8NnZCCZMrlK
cKi45d7w0OloOB7CQpHM19kp0oQp8xdoZ49KgMz5EVcIo9Q6K/dwmOv84u2/LY8E
x9Q9nBLhw4tOnLYdGhN/c+mix1V+n8Llwfr05lxYGn+cr98LL/En4Bq5v+AuneEL
4/fxLXHQhgoXbYW/z6OrepZPthlUIXIYXbJMle5Nu41RaEm/cxjfvUPQVA3l7y6z
n1cT3oxB/ozu45nfZaCl728hGlOueUbf+bYcaC63c7Ui2OiAVdgnoszbO1fHXVzV
Fy7Teab5ZS9j2IDEX1MF5i90C3t429uYRV3i3VpDmpFDoSq+oGyGq7KThNKEqIgO
l2MXfxrsIIrh3V+h+Qm2ycHTGT02zT6HZa36hlS+G0hi8+tXIis45KGHilrMEbqM
WFkaOZE8Equz5UebMzajTaSePUyLcLT5qRhizhJpeSDb6bo+uNnrCLEcLvI319/0
bMuDZujDez5dx3auk9AsCnuEb0/5fNzftZZoJwjTyl5tE1KwiDAauW5+Ohv+Bngj
CZUeI4VapaFrQak6cf7XJWWeCD8iOa7ALZnPa8ll9MaW3N7Q9vfcUI7Vv2IIt5lr
hXASkNZEZPFDR25aWCN2bLgv8FWbV2bjxYRg2kbq5F+cw3weprSR2j+dHAzQE/H4
c3UmgTIjO71wjiocNmKxTFCP4kQ5QDkLoXBUMea4g+deKbx5dEBcoN7zaZXRUKyf
SNb2PEo1EdRFHjSOpYdZzI2JbN+9381413IdQw9n3y727t4I+MV9jNMd3pReCXWY
3E+tguE9UTXFJDa5/bJYJ6pjxwhxgvaRWxZxp46fzPm6osL0uCcP7sngy5x0DOsC
E1SECmSoJKw6cgNxb23kon1QnQF5g8rhbcOnaRD2huLATmRnzEAvjLjyXJxbUvZo
GU9pvkbGSL8lGq/4H4qNJgzhrAygU2so1KHAyxtO/114dcz+HFgehK4438bcOoIT
BWRZ+yML30LXDNfF4neKDrVb0WiHAYfpjxK7x/feE9cHY9uoFhZArsBnfTybliwP
HADg+5bSuP+l9OSe7n42S+ejDPvj40s8AV77pnTXPkjUNKm1zUUKAWnrCEan1OGw
2CNpZKj2rGQ6Vsg1hycIHj3gANy5qvzF10LQUurcptypWWVIgBP/ot+pk2Q1k31e
dEKbMGOC5YqSZWteVH7VyXHbVT0Gq5JUkLc6TB4lhdogbynvbKFAi3OBh7RCwBys
kStr4Ia3PAbKefscQm/Yr+6IhMqJqtDXTgp/tYC5Yg5GrDjkqkOWIIsb9cTjazFV
UgoMzre3RtYpNneJPkyhVYaoZPu3eWz92L9W7HRfRR3riSVNyskXwiLSFDLW99ZP
U6OwzfoZiDpQ83sf/pdt5uP9+Hf4Jhms8VQdgF07EeEtVyMQJcEf2EQrFw6bhI8R
ATCxOKODNdBQ9nOvtXFB12ctgSB7xUswxWsLeVViaSIhcTPwsU4Bw8QRLpcP005U
BdjKCHhLJ3lB5j+8XvP8fiSa1TVXW19gPYUqa4JBF+x5CPYAYxpK+WRhkem/UEvt
YNUj5O75/1BGRNpKsdSFLPbumT/0IODgP/P3pICaZEnG734Mww+qqF9sHdI1ZC6Q
jW8J+Isg9ou/JNY5ka/toNX/0lYMyCWWi/9xAVnYp23LtGFPpxVKU7Il+u483QKR
H6YbNiJWqobO5zUv3Iq5lvjNo2e+FRzrlfTRgJo4LI22LDv2XaivHuGJ/16ZhLq/
a25LGQHzzZnC3kqd3A0S2oBz09vQvQ2Srt8BJF1MbOl1Z+ZhGofrC6oIlfHxGLk3
oE2GJFlMa0QJ7VMohSKUYbJU1afBRzPp66dnedG7TXtk+NvGCiruGmq4jmvw2bYq
ZGe6y1VoxTtTbyDGfNFU4OTflG744NoCQGPBJiur4OBXubP3xtvnxiRNloXi/t2m
PfZTNKt3imiyAHuGW6xWI3DiuYS8mHcvcLPH1qeY0I9eidGF1NrWgteMPP3fksfK
juZCxBY5FbtxuBtQ85ShbI3Dhd5f/3/QOmozuzW5oMPB3agStqE34EZX2Ms9dey3
Bkb2QaKQixB3ghzmUZA6fWhL/uUNhqVVl2grBlFZZJr0CoUgL6s8lZIGgFqLOdSC
1C+//K0WB80OzpF3kM9F8QFiybJseL4OmIpQwem3pSWsymWKK7efIHi3NbEA1Gpq
LH6E44dStOj99OiN2u4SI/pAzaIkCaO6fTnoDCw41shTpNDTid0g1x8SM7b9pe0O
RQQpotHDGh6AqdJ3BWHiU5HTyIIa8mgLJ6+anoGV6UQXQruc4igXPYZgfXODMvYV
8FDgO2urxrdv/dYWVIn/YMwogNriYGd0R4XsjndkEcQ7eaPeahbwGATK72xaMXTl
qkilxwAKR0ELw02tDRoKXBacS+JG3xpTu+SE/awMrlSH/t0bZsFW/4fjQ55mA9g7
HUh6+nTzs5jtI5EqR2QXHNXAB56lNYTSL1RIrCaboW3cVk2gg7CEJcLZTyVmAQd3
wkc07JLjuGelnBH3gLlPyRDXrTinSZAlbt3bz2hrTHZd1M0cYUFgFvZdpSshpo3W
VJXLJWiP2n0oPxkSulC5Y0aKlx9UJxfyiD5/54vd8104EEHCQine/qooYC648PrM
ZPb+OsWQc4zfB5GTpBNMqMJ6teyscLt9ZCVZ9Lu4DvVGHQm4HopWubLpM2qk37DS
ZSv+YNw2f3r6c5RW8a3zs8+mERPEHe2D3OaYf+WV0kgy3eA2Y4z/XwlgkTelEyD2
tdJz4+839nzm6MVg4fSBwWmZN5pTW3IhcmPjnBn/7u0F3D3Wdi11YXe2o23ik0fw
IMMTjmBlvLWToLNvy6shRqO7tBG9QKlIpKi2g1NKcokzeSbpGHdAELw7FNyMhOMq
ELElYwlLVJoA1cmyMwHiU5fOQBSNPQ/hM2f2yPdxWxeGVGb15C9xRoHR4O2CuAKF
1eIMYWrtWjFwXd0H+O15wBVYMnsuv1RGL5cMNHWBfiIlIclKEx9+3H6zbN7++Ewr
VTAktBTbwWgF3teEnNV4kY3TtXTgqCsErId9ssCbvX0j0hBOqKujmfXHlJizBx07
gKhWvd6mvBSRJNZWbZ/viO7wAoLyG92jUG0enuqGAwlUIeqslQ7kRI2TSj6zy8mD
bZNrWDHWIgidCxSTi7B0e19dZZB4daKZK4Wh+N0P13R5TwarRGL5I2IszYdFab/P
Oem94J9VCFtGKCgv1ZL8SC85q+NW15YCBeS3QUspk+sHrslJzVzjkVGLPUHVaulr
m/Kc7KXn/oPp9EZTFHNshAG/b+9i1GISbH+7U3QBNxh4siSQv9hC1X7DPGCelOZo
KN5WAVlxfzLOJiT8hGbZr6UleUuXfcBm18ceCXXUZ5EY+YXzbRgbBWY1W7Mt/LGh
l8hl84+mpC9xR/10NhluaReqsgKf9PfhWfsihK/w3C9IkOHpc2zzNGFl49VYp4DH
SIwJYJku4Zs5kzqqTuo1uFuoHORlCP0ZMRbUCZa5Ghgje9K7/SEd1sX/aT/soblA
a0ZaIhxVeZMXnA6VPrNqn+VQTRAItMnSflEdIu9Z7AM4r7ooBNHnFSG6UV42x/Ze
Cl59TKxoo1doojT37v29GW2gp8lFmvwyikr4U56Ie1W88p0MNT7P7/nQwNHf+XPx
zvAPJPlYeFwt3VITprq6CQhRAMzCOk+irNyHQg4HavBrWh+pZbEFfwWNoZzff4UH
/9trM2YpBuHFsCzwpDf/hk3pyV8RTBBCNZynzes20gdkuMpqnnwPOQIUKtQNE5Ii
WoTu60Z4GTZuqYNWz9eqH8jfdo8Xc7A210Oxax1V+JFNDsdIEUDkaBLWihG//HUB
Ao/LJ+rlAhED9L7O2Y5U2Q4a1kzBw2ARWlkbY2yCi8T+NiCLpQznCcIwDYicmkn9
8j6yX84Zie6lGmJF9lYXIgGovFcIhFlVZDoxWwtJzJ7D1vfoidZ6JGfXHfpZOKxP
NMKuzOktjBOP+BNblhwTrnh5EUDXIqXaLXjmZopgtdNB6Ise0fUPyHFFyfiEfL7F
UZ8jj03gx8/nG4OGsAkZsk2KoLtGpqAWRL4KfYbgdojya3Oh2jCcjn8/agJ4Uu4U
bOys1k1ceHXNmkSNdRbn8/jjmQESomhTxwpuc4AHj6+XQFoPTB7gcBtbslLgYouG
qbMHqrlJcNHZaSt66sE0RFE0P6iTgj5JlBu7EcpNr//gRNM5m1YWJ1iL/zxC3h/Q
glZB6z6x/vlmWhrJX8OOa6X/ZuJilRhhXJ14r72rWYsjQDW6KGxCA/hvgG6DXJbk
9w/AOgOFQ3MfwyxT7BV1H0tP5AGCtrC9NwtU84lKPlGlENuYpqH6qj29bI+3bvmb
yatmF0jFCt0Z4GlngrmHf0F2KFRVN0QyZ1HOwBnPcDCho7M+yr6YJwrha4jXQLwM
pLDY/Tq2ZDCY8yOZd2J6n3AN1MvSLwy43yisAxGN0Z4wWLmVBEpyaYXfaeGIE3sA
CjxbTKWQ1mQSI8alX5/j8ES7/+YFaELNWp/jGc60BqtQg2r70f5xkIe6oa8nGTqy
SfkruVMq9lMJTOoLUq9XPr9DgQgxvbf6PgeI4usEdNKWFIqy6K3nI7OYq5Nw2bdy
quRXExXlc+wBTCqVwYlBG81uopLOqzk/IWJdhMlgocBo7iMySGjrd9j7CxRJ+N/A
6CPw9woDPKx9h8jEDQZeafxtsf5IT90w4bOicB8q52Ps3SuVU/eJH7a3PVOg/KQ0
33VSH78SzNceMR9waHnjbka4KRI2OVzoUS0wCVMmcn78Ykm2LvWy2KYlMLGdZVtO
0KIO5UmNmfdZ9flYXbDAn9d9pBm2BMkAWHVlSaod7qP40/LNlr9KzJS57ZxHAb7P
qLjFiF3IXkH7PDLGa5Ge69ivYTMqqZlHkHAzlrzdSAiRwNK9Eql4xWo6R8jFJ6jP
r9DiG89lO1qCz1ONBM3qlneZGwtoSzcXmLJrR+bYLJZhWgY/BuN79kpJj+uXXcYi
sXONgQwdRqfqvEePnLfU4QvXKM6E7CDdOdu4JIR5Qvq9uSqQdiVAdHw+n3NEkXWJ
vXz3BZlYG4sd40Dx7XKMXkXMqjv/ec54LNNdR3Nl9iqJC5Pem9RNYoXSY9ODVP3r
5I4gP8VjIyO8zbJvVYzL2elB3j58xDsvkApbCdxMPHf0sVbbpW+1/wA4xiCz6mmM
C9Jh4JpaEJzNj/tI7N4tRKu5n8g6I3jhOG3EUijq1J5gTA4I7BsV8Sn+p1NelaHf
725kcrOlH+z7wi8TSDhahSFmVlrrEpXh/zzrtaZwrXtWyI9aAaGNj4kgjs+AZvO0
/zC5I8hpNd3r+Ns2p4mmsJVBq7WDbU2zb2WiX8xOy8iD0PQmBEbmi297I5dcO7Gu
lMDui/BOkKTNSO8inklIj1YdTtcPoAfsBh0WrxFrN2hEPo1sGHBIhCo9ZBlSh/s0
aqu0W3IlxujkjPQe9fEacVC5+EqrtoAqTOiHPxyfCY5QKMQsMv0DDUhZ8IVMuVzy
AuXQgES/3ropYBlljMwjdKyT8tWR8oTM4dygAW2ZJ3zxVaqdnHTIBAxNwjVDa0S/
IOrklu1BlQ0/uCEa3VvynUHYZ9fIC6iUBDJKslYPMGpx2sef0sboxyi6akaUV9ZA
HJgJJpwskwINwPr5ZXc7a7KSi6PLTG4MIaJiYEOxX2YFFYytZrk0ZBMF/WhYTSuM
PgR7HWxhJRaXSa6P0leI/vopsA7pa28E+tpkO/Q1X02VjcZWoyPVP9PJzFwhTF//
VdJbmwbrAsrklYF/mtTWezidSfd8vDMEFPb2suupxG8ZeiaEn3Tz1vZ35eLwzNJJ
23JvuBIH6s+UuDVfl3FeKsCFA+577Cg4+Peq5obxG9ATFY5m3K92TjGDVU3v/32E
JrbdE51GPwrDDjzspGDi89Uwips2/ILnXKp+xhn1kNIGKjhO9TuYwUTkpkzSk/j+
8X9IT1koKD3q4pTyLWaS1jrvlo5XA8H90DvE3oWx2jnHvdipxhUT+Kqjrl3y9Yjp
ZQr7yuK97niQFtZQov+NqwxgdWH3zorpALsabgUYIDmkc+BZ9sYM/6g6nxH4ybmR
K+pHldqFOmc80311az3IH4ckQXUfMRgZNIJ+jrOdLOKl6SCODMC4GYY16RclyLLl
0BBaQuqAQQ3Bi5ABcQt4QR5xnORGve+zpiggHxf0CZAebyY7SRu4vqmG3I0J/Cbx
7W46KPCvWHUDiQBdT1IC2kQma8msJxBoopK6Cd3je8LVxmyIbuY7zyAF4tXVLb4Z
j1qysUY0CxyAWvg0gV/KZ5/unu4Sned62z1HmtaxOUpz3LCLdEgbQZH80yhHr+n6
iDsYSccu/CrxoH9C1XXQ2MHOAZbPY6sJ85wAKQMvuYrpOUhMqjswtZnCbdo0tOMG
d1xYQSY4dTUlYx8zlwzty8x2Qphq7ceECya0JYHJborroa971OwQZMXuzQlofjz4
2vb1nNAJLUGbsw3f129bMUcBlG7tQqXqADAB4w1Iim0VIZglOdiKEwsxzRpoVBro
feK93tPMP472GJpwv2KN6la+e+TG7O5IVXCEHA2B16mN7+QRL3NGT7nCaMBT9TMQ
JJm4Kpwjl4Bq2bCjsrJM5Aqsc1Ff5uDjvhBGOJ91gopUTSnBK+DHMg6l7jkNLDdj
wHTA4wYfbZrWig3y6Lnq0Rk4/DGuBlvPAodwdwH1bATanf6afPYv8A/Cjrj7gmey
A1EdeZKylcc2hMS3PIEtadljWwDjmgGfMVd0qAEZ0yd+uDX70Kyu/GADHHVpXOg4
sEDYn6XDE+N6PoID4fGHcpMZ8vNbaIEd68ZvGfySpEmfO2ZK0y1jI5e91QKXFuTs
6J9AlrBKbcTC2OOwNRVbt//0Ada8EACD3MwaXrow1Hh/pl0bCqR3jQXUcon0iWq6
bGSczxh3Xn53vy8yd/BSiOs99s5oN+HuXOluLIqlitbhYOFLCXWSWhbJPWNuM5Al
ZbMm9f4xDz2NxYRzpMfPUp5YIjiq9U9DivWJib/w7Ci2JO6k5nbyUJXQAgXjsZIf
B5xTZ1LFhQduO5QBtEizwWNHd65HX+Kl5+/yB3NClTzoaL3almB6VoxAyf2jdXPi
XTW0Oy/iBhKBmzshZLRtRXd7rBSn31PjgxcWDb5Ek5NwHznZIAD2NZgkH1Ojly+z
`pragma protect end_protected
