// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
hGKunfWVBiEX1eQE/ZdaLYEylg50W8k8u/ag/3iL/wXGwr/W5tlQWCy2jG2OLRjCgxw0HQXOKNlH
/nKmnhJ/3vt7Ll207gNBGRcB5znSeTsnRLP1Cbogk1ooEb2Hc3pWGWM4QJ1FXkkI99rY3D77gn1k
yYIyVXDr/DCkunb/RaCvyxYddaCqYGxabElFfGYkgOaipmvr/HZiN4nLvwjihDnuoyWmE/Nfqi2l
uEA6FS6i97LsJ0LIVPPSJc57WxHgsAEQ/b+wPCHitwt+HNDDJGf8rzeWCRRgehsmtkn/nUqm+5jc
OGIqiHhKIIx9odYNNyCNrK1M6PO6Tg9erPwYkQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 25104)
sl7tP4GkCXFKZurMHvwCwasZNBRj9hlFrqX+HnjRYpG8fJk/a9wz5mGznvxWWzillSdQ48dKT8gN
4mO1b9flSGLfu77RC47VssYaNLoIwghLps173XAnZUG/Uxl/Vo1XtABjpUdsVu4i8ziVbCzh9IPQ
EmMM6u3B3mtWMqZqPni6c62VClHIlV/xO1yOpZqwTEZTO6QYLjuumkenxNcjkFhVzOKuSSIQfM+f
boixou7e9y0d5ROH947OnvvClFGf0PeHybRp9O/CmrRFOMKfWrH656TuHS9QClmALZjbVUk8aIHD
g7rvfL9RLTmO38Zhe+axBsEWlzTDnBFwtdvswrbt+LOZstRaWioCov0E9lG1p+cPGuQY/Fm0nlrO
La6+CGTrbQb8kGu9pB8x3I1TX2qofZAcCA+VRP64qhhydLWL4Ms8vtVOMXiRpZ6vDuQ3ZgMbT/J3
KxZBisNMqB2Sd2yoK/WMpvATR8n2omn+qIC4qeC5bGhkFwUxtOpAxAEGrSE0dPR21Tdgs9Qm3fNZ
6cGswizx+PcbEzpgkinfq5DwYQaVnA5qp+1v5qNOdJQsnSDJILMIp+XO6ZLW0pH9B6CcqBwEvFUQ
DHu70uZd71ItZ7Ii09Qi2hbSUxG3VofP6sK8ckoCvnpBHFNNaUHi2feI1PXJIugYWetLE9sx3DQi
5+RFy0vfupCEBj9a3Dq7UOew0A7BJANEwojAFV1W+z67q3cf1B77VRep2hYi60crd3UeK+NXykus
6fCxaSunuzy+CX11975svuASvbR2GKFOt7uLQie9tyQaqqk841fY0W5oHpZqkMlQBDgHbXMhM35T
hTyyNx0PgHIpbR61seYeFGvWW6fIkUmMdkx70mUL7weWF9uw09FwbWGrPWNrFQofDH+/IzZvnGE7
P5yOGDYzLdyu72rIYXh37VNUmDqjftNIr20Sk13S0lYCC5VL8shZA/XhX8XhQyBY+QtmgahsgRzS
T9FC/dFzfIIPsEy/WzwmoV3+SYX7csU2IpEwIRoPVt9TcagFz6R8FUPQ0sw73Fxn/px3fxrOfs6G
qVF/Qzo+WdZuMPIi4ZnkiMkg9CSXtsn6WO3t5iwTzLdD9rBMy6CuH98F4Y9XFW0u2SAM3V6BULaM
RqSdGdhdf5uWmWSlQS7pQPsBprmKCouqeFM0/hHB/AzA/Yh1hXAAwpJLuj/eC7BdoHGbt6/2nlBg
7/65Ad5SFNkYcpRTH+7RT4+IuF9NtVoi9wajwYwOckFCk+QFwCBi7Lm80S+roXiaw0xjcNissCLo
AjpyCFcIvV2kB+mWgijWl2JbKdrToDarqp+jYINF4VTKj22hkqc1BjeLhnJmXybT3cuD9tVkaUKO
Vd+AK7Yiv8EdQQWFjZi+jpTxjaerAP9iTUqwelJSK6D2iTOkRGUujZYeAxK8wZOPB0Cy4klWm3LJ
0/4IQFfAkSPrJ2R3KelIofuMEEaIlB5hyw/sdWhznh5XH+rHgdZsPeOnxctoKiq1r3eATrJlnMfa
jbn2eMHjrYV7TV3Gpu06DjH4GhTpIom+87xZyauviV4ZPVuYIjQ12l/3cckfGIEbv8moVyY7VIoc
xLdNtCoh4yXU907UtIA2hnLMLWK464iTRZKGa0PoyzGNICutjZElI/jd85BTA6u7+aXMzhSmCI1J
89fJfnw5uETkBsKe6L+rb0JmfQa1l2NNIqRYMGp8Iib7VoTkw6cSqf9lyFWiEp/8YEAYJmjKwxdy
eWLtSmpGJfl6dPX4UE+x2l5ZpwPcKsrZDZCOT4ho1mEd4yYja5nXLUxiTk8omzIm1z4r0+zpcWy4
R3DVYGJiL7rH79FHSvmanOLKmPdg9u2ec59yzkZERCQ+oXxFwF7ydFSIEysgAHqvvDttNM/k2u65
06vffRbZXxUG4gzq0v2Gq+tgNpBofZTyblfKryA9FBal7JkNkRI/Z6Zn+W6TBCFrXHOVsgHVn3ZM
ClPZCUNTSv6rhbvxdwD7WMP9xmWsfP+i4a+SZP/REEafQbwNL2aS7oj2W8ZsAgml3u2T/74GrXaN
Cv5tpLLzk22zreSFE4EdqDjxGUetlB4MK/W7AeJOZZwveQx9W/u7VQNR0qUEyCG87dXizTavqNtW
X38nq4zmzcpYXRNef0KWmZkaY/3MY6zI+6/I4K4O/WAJ31KMs82EO27fVRboHou+25zYD031zyET
NNN/jVdLOkRFEaWFXiHKrwMUeE+acZj2vgX17sFNErzpbhmxFAHB4DDHOcmzDpKARbRX1kfQ3rI7
05w5P4NQvucJLRhWDFXavi8Kvku92Xkhcg0N/YT8uN1vsXCelCtiExI0+VWtiZxeoLFR6+Et/M2t
ub/SEqE0fi/ql6kdmW9epBocTa775hBPJh7UugWu4OHjGKvyD7EmRif2O7sgQDU8MrtCFGdO9GG3
xYXFDJtLl6WE5u3Kjuudq4FJerT2wLscPApsmrmB9a7NrFZ58A1YCuuSHMW5Yw8sSWwNOIRsaFCE
0WIiz6GahwGBRMJBHwB+JMSXGcLOVEtBlYcIYl6+QMrj9iEClrCTnKJlqioQb3re2kruIwfa0DeH
hIXxaT6PyzVKr1y1M1+awCXmhySX6lsyOWMpnv2fUeilRD4awlUmXZ/Pk+0E9qr3grMtsvI3V/XE
UIfkZNyKDIVXb+D6ijk8s78cRTSPj/gV5VnEJEPDDKOT5RE9eSTCj7PaCKtyQ2059mRBTa9XpFTi
M8TsmttjfPuREVJcRmSzaByyVQzDlw2zUb5TlJPjrq7ru6wOELsgw1ZGuW8dhVkJunQ/cYjI/PWT
QQ/TFMNgnEiGiz0WIjxExQb/CDeSTb1vYblejEWL4KFBEAEFB1qEAoe9Ivdchrs/Ly+C79kcYPo1
sQczz7NQbDA5j0trA0BSSfQVCnghnlNX24nhf0ydhYnddK/b7lehFUTODckIZxtTf+PVYjebmX7v
SCmHnRI9aA5YFkISFtCvaTJSS0GwtDY1UMJBb3co+VC7MnMrW/eF1MQMSRn50LZZ9pVROPlIy5Gi
nYNVBtD56awltY9olOZ1poNsLEnKBs9G1BJypywU6cywAeeSiR4etHHkkc3+bF70Z3NMSQGGNzEQ
PbpAj59XWFLivGMA1f+OU440CuScFimI0I0wAWJKk/HUiI7P8hN1gygN5jzNJFK7TmtfdJgBgjde
+CpXxkAXCoSIVwcPasU0GBiq5cbJ1VqetyEDrJYrHBDsnOrkUQCxkR8sGz9mClEuILubcISs0G3Y
1gOin1YzcZWOtSFMsv5FjUscmb9TCIhWrKLEPq5iKiYvYy69/Xmcr+kbWs7S8+3kop2zgXQpOnzI
LqtQPC3zRsuylHHivjjuE7PMD+BwpXgehCkDsd9orxoaxQUeg6mt9//XoBFsgF8iPUm0PaZppH+M
OTvnPeYsLCzdkzEDM4Im+EpU39s+YCAYGoD+ZRvQ59STFOLDASIZ5mj2Et0sdxSKobSamjc0D55y
jFCtopyOb46TBgbbKiuSwA1dUj+v/JGwdrFQ5ZfCcW+ehK2DjbNsqa71Pg/lYQ/RuS/zX5jzp7+H
Gj3I+vHWTwYfgwMyyEyGP/Kd+ty1Hcv/5raxbvaBW+0FMIdmRvteIDfc+LPmWYfauEUf/dQpcseK
UQfmv0L/wd7cy9gioPxf0QEE958BcTg28+ZeBWGksTAgXKVmt+LfaLqJK8MpCjv8mAyCF1JXX/zR
hFQ0sGOLW3a2Y0C8Qk+hZHCk3E8K3dhx2O6DWHH0l7piqLpxu9GrlsuocT6ppYUsZGaiFTzVtzmF
2HWwInkUdu6EcvxgWPVPTBO2eITrBph76zUC7oFWMIzjUinJbt3CskP8gHj6zkSU+DDlT0lXUoNe
Unhaxjd64GCL/h1DfZIV8wrkaL2l5FL+1Spa0IfNP/3M0aOOr4/sFQLmtXZWH73G6P/We8TIansi
egjG1chJ326+KP5PHQxU6ESUlanNRxNxtdvXu/HcWqoAPJx+9zciDYR72N0WZnCZud0oPPhP2Nxe
26lZWLcGtXI++bwZ+rpZseMWuoLgmUo4hHzqfNlAMo05FFAVTb/kOss7M7Cr6y7/EDjDazfVWVu2
AZ3bI9Q0I1nMjXGnmlabA0QsGYDo1MwwwrhdKUCgG3jgEzPRa1rEVWS66HcJujZ1/7QKoDn13e8H
N+Fj94OoAc6+9Jy/alJ39ZVRk5NNmVr9hZT4ioldV6CG/AsaCvLWjif/m2VhAV0Jzp1LwaiFyULg
ojHaUnCbRHIUhqaS81cDOsmi0c51tSEs5VmpZCuvrABkj5u5fWYpZiMGjTs/8uegyrSRvlqMxY9o
oqg+URrXLC8LYNjnHPEDPW4EcjBVlSLUnx16EXgjdWY9c+MyxSlo3RkOdr5oZAzroz3fA9MsJQs4
aO2Ka4NsnDuZ+rkas8bGu1UXHj6CK2NKMUDV6upEUoq/Riy/SbN2QkOufFyrONPrZkdM8jMTuJmX
SB9kmbWYP1d2d+BaO9WUrUyTYDA+zw3/P224aW7HqwTohXQXlEsAwMTQg1TtNxVznmYyAF7gt/ty
Cork2OWlFLpZEhhxV452RL77DwBntkQq3TE0th1kiYmyn3LHZG9JDwRqm+uigWNeS9wchxTmFfYg
nQE6msVXTSNJnGFXJulPnKTui+x7VQxxMmA951bvFrcfnXYwvGt8nztLSOdDmDncXb74vL/j+3NV
4nYhfKuVKE27I2sMQiR3SrPZkT2W+YT1PIQLhSHpYMHt7lzTpNGzvcioQHq3PhqwLG0/LQncLaI3
EAP8aZ4AWbumLhpKkxGlaaWgOl0ujbmosBC3tp6Mm5WXNO3lQ6VSwAXFjU0AnDpYWDRiM1cFxEvR
MurSfb+eZgLmBplOc3ka4hSJ6nJZ6++HJhH2SC8vtlKx4MWgM5yF3XLvXRpfEg52Ftb33GG579lW
HHWLH7xymZ8zV1wkMcqd+ov4AFYKTcZF22mlDzwnXKsub6JuqLcxO2vbVzdw92d5nLk1cPPnOFOh
kWDlw2HfFTv7xaRPBJIdmlO3gF1cNt2FCt21GGkKoQkMrljiFuNzkeTmqG0qat3fYvDKcfSpgBgP
HqPbqUEfh38yVDtHGSRSu+OechKp3s8Eb7XzzqSPiejLRXjcMtLApBPNrcD+oCqRbiKUtKanvK4i
UI2LKR4cJOd+WGxExivu50NeTI70CxmGOpa6dJANUbsci4s4Cb4YDS5DA2fQ9pxmm0RpOrx41GyK
6CT4Bvl8EmnMo5TIcTENhsehkJ0EszbhgP53/E95couDJNDml/FrIl2cILGZlLrNzsEI/SQawp3N
L8jeBnSFFABo2tpLvNEk0Ynd5rp8Ttmet8aNhvo2J/LrzCGVXdpRa5fehnk0eMw3JOPewAJkXaB1
Yrn73fcDUlBVvaVS+0/5q+Mp8fKtF0rZDXtL1T9Owur7bszJJPd97G5S274uZNJZ4+O3WVmnscrT
xIMiJakemsN44mV6NFLTGiSKFFgQf4SVs5nT7QGSObLTZKMWlufzekQoCRapp7j0URRUY59xqsl0
OazbOWijJaQPvUOSG9rET4j3+q419arcj9j6ye10nae9dOrxXzI9xLHw/z8cqqBaNco8xxZuoOPF
lLQRV+aIs4qjEbpVZ1V5TuKSBVx1Z4vlAGqk8M9hq9jE69iFuV7aMqgPlomzziApE91ugdGXXTSJ
boftA1iDVZSeh03JB0iiTMKk/Y6rTpEqwaGKRDlcpZmmlAZ78X7CBcnnVyfFXU5plHjle/fEf91Q
esaLA2QwgC51CtC1u9tmqk8Ejg8PrGySEGxSQSU3nmMeQR2o7oXMOXvsCMJ0/+PZMNrxesPd1cGx
OiVFTbw1vnpSg5C3mNPEb6sFASCdqyFTcoWTe6h4j31S4uOBxMxBTnKnaOfKem9Fptmm3ic9tf58
yQvcB5tlqk5rU/FdSCtL5QEKKia/g6W1gC2rUrS1+fW6Hz8LlwrRwgLVT85w5NDSCT55V0jI+5zG
gzedr31eVaEBV6HwEa4Wj2z1cslRpIAYC4Bmf6/KDQiIUpacumYOwTNYEAMfeimGpYq5aHZQNNTr
LGrWJdFaNRqmMApidqKT4uSRwT5eRVRkJzL5/ct5+JrBvaOFmPHm0wffgGlLW+gt3WknGG+hn4so
i9pOwOZS8x9E7AmIY0yy48bB0Cku/w/6AAUS3Wm4gh845gpiE+mkgRyQr/I4j2Z5JuOR7CEYziNz
cauWJYFjlnaAe8N+dX4w+FpNJiYD7ArWqTx4ET3LkavNczvQJLbEJo9GQbZPpOe1/uhM4iiCmuTU
KxWVBGaOoO6IMN8CsOZnnb+UPx9rKrKYqGrkLVVEbYJX1Dg0ZRvj7leNEbgPVaHJnlMlaA+1JsrH
s5u8uTBy+xdIbQcstN29E7DWnkTHwax5aZiZwlCgX0eVc3IrBLvNicKSld8x/z2YmeyclrlzuhFV
bM3CXGsp/mhqbeUvEEzzMRj0wwUj3p1/8us/jbIBloP969I98k/4jgO6At/Z42KhRfQIthIWvjgn
c0oU+62KfIdEkOGMs5wpK8dwX5K1g25+wApzSWUorPlfHDRMiEh8xeYhJgEWn3osIR1/nUKBp3De
a+T3YxamClBuHy4BywlC0dohnzntxj8UEU9E1pcCOWDWp+TNCPgdQdK9XuZTV98AGbT/cb45yfBq
Upbe85AlM1GmGSb3q7vmc/39uoWbH+3bpFZAp09HstlaxF2o1OnEw6ONHEqM1elO5fnEVaUeOFXT
qLveHiUAmkUTQw49TaSgtz+G0oE921cTr/WUb3v1r8pi3cYRH0GCK/HL2u91pe/tN/zJUOM5A+Kv
9kL7wGc2CojF5NpFnVRaMSZn9Vu0EFdd75+pbQoPkJYAqCZ+dY2yaK7R45j3tR9QbJS4ZZoZvnOm
bwheCS1Xv1el6E2ET6l/bLtnxbxXAmLRlWpOAAVAz9WKL3GGxWoM3EzB6PPea7F5ehLimnPADUxi
Hik37GMYO2RXTBFI9ZiIunBv2bjjthBZWcmqbqtUZIQbdSzjnDrxTxKB4EPVd9j0/q7QPlqbzhYV
jnh5ITMs3EUrDY5Gr0GOB0/lQlBHlLVrHcHW7wxeDjOHZz0iMpJOPEEz56GESILi3nyaQQ+RQxNN
71ljM0K6Lld3FxZ7BGF/qENBSXRw82fnoekWkGbZNvcCmkAkI90tjJ/LR8UjXAUWBnT0wEgnCs0O
pQp1aIuZtlxXJwtzlUCzdqxHXp4aigIToBNu2dQzlqB3LuiBiflOI98PbOm5InDrRy74R5wWeHfp
DN3KLfGYANJA2Qx4q/MVmG80PzAi0Xh7HhNdVzLtGpyfU2zhEqcjkADejN7HfccKWh/X0c2vVWir
ROkqCdHdbYw1u3MdhClm80FmLZA4H9KOy59RMz7V03H8CvFhTcbqlFfW1Sej5ioS72TJyf+vCZYW
WqE4MOihBnDXEfiY9BnfsnnfbJ1rCKjvmSX7btsR5q7s29oULvR2j7MGKeslNXg4IjxbQXdarr/C
cavwTybJm7akk9BjKWHAupp+Xhq3w0NYd9nHMZ61UGA7LXfQhKt0xT0yBYmGZDqe8358xvXHnB4R
9CUv8X/0pzqxxz8Bpirgx9md1Z8ix0dNqun5P4ChN0ojdC2k81QEPcWcecQcsHZrzrT3g0j3BvsA
bDeoAzh67HG82xGmhuU+uuRDF56IlUkwGcEZz2w3Fskk60kt53VmNKvj6CAF+4CYhIbsDhWOdQAg
MthoS27mix3yXWo+tyTBBHZ6usD/JuOsjgqFM83BIg/NQzp9qDbAW6VJb8AXd2MwMPczuIm4kP8M
H0gmVAPUwY2nkVSY7y4jJ/xcYzDd2DDfNr17/nqk7KoaweIxuZ/7MasYJgWR5b1/cnNQUQiBhdi0
gt5N+e/2AfS1RcRr5Ebn6VXddK1Urkw+/ePMjyEV79ZW36XT1S2A8oMQJRMYZs4c4IlaqWwhuFWa
1ih66KEwLG5nb0OtGGRJTzgvO1aDkaKyqArJ77sBCnRsTHm0GTAX2fzWvyCN0e7LddNHwTGYgJYQ
mWXY58itwzKYhjxf82u8JWk8892w5vDTA3DMoEuBNNS71ZSK1fRrETzLQPVwAXHcKSwle2QpNajp
nI8912yv2SM+YblpoS+SOksLmmE1mikvD/GloObcaq1ca9x2zAQ39P6JtmqwyWlZTWlU1s7FEdUf
+oJopPicMbALaWVDLgMTUS9vWpCBJuOG/T9vFNFrKAGUuWjWzIh3tjkjzgl/fKW+9Qtca3y/fPyt
jGyFjRNZ972krx8wgVOQ7drdm2ZNHnYT+ouVb8HlhBVdHu63WX8FoZ870jN/cMhUykwOH6XG6Djo
Lc/iHVvSSkDEH0g6d2KJkAolCFd+N3ZdrzSpqsyXwRS095RKDvo3s62K2a6Us4F3ekLY0Tl6huQm
5MHrJWbTTFdfrT6m1rxkrpDobt6QDof5KRY2iOL9SqqkbxZGdtM7aCIUDB8+cBc6LfqM0jF8dnw2
gR1HBufJt0hW7GP0PVppU19PKw+kmUj0vGd68/wy8HnjKk3t4v0ZdHQoNnQ+ACi2YYiqpOYy/P+o
ba/hGJm0xGHrTB2HTVgH594HG3j379FsBOsipELcpHSty3AHpgEAvXaOLBHmc2cQCg6HPTWM6CmM
rrGHOkkljf9Ha0VnQWGUKO2uBc74Bco7da/Qj1nLcKcgzfgoiIdwdiFsR9/1SRtp/w1C+Eccqlnw
xlhbC+7OMz1Agy8dU4sWAETBuZiy8j8y4x1i10Jg/Uzcbm9oswg6BqXUmFlRhfkORAwo12sihv0U
iw6aJ/dtTjPIh2yTZSXCpbHgHoq3QOgNZZLOj76UKfcZQDYZ7P+96HErmpu5lVSP/NlcxAzLnsEl
Xt/+Ee3kvLQxF1sPOwu9cQztwqzT7E++whOk5bZPwc0GlfZ9j3o6aRPPyM5OiWkWOSUYwN4noilL
5zKLH7pzdczqGgvjWFsCc+02TnxgabWeOTTYYI7cOYOtNcNps5YDkLYJA9ZMFY26WP3qtJ9tRWzr
HmnsP32fn0j0iFKky4CNXAzGl14trN/9tDmSz0ud5yWNiwDPNVDEIGlqTVX1xKGpUqPJPLJnqkBZ
SF50NVG29tbPwebm0YurPgTkPa5H91x8UFaR/mYT6UfVp2nt4FXILU8tZfwernY78avF5ZKgJ6pB
MDYPVz1v9S3aRyQ0v6YBrxjgXi/I4M1/znu2aL7WbF/FPCR6WWajtXEnE0XSNnvXRo9WwxqlYNjq
Ke2Q8s8VKC8pTkYKFvvYdNieGIRUXx9axybFB3OMBPwy8jXksj13Gdhr6zXymhhjGggbzkgp0m1c
wLjW2sJj3VZgEsPcqIscDEvNlTNlnPwQcNM+OD4k/iUoENMM7+f5TQkIQm7WwiI80BxDHqrZckfl
1TUMwYQVW8jXkYylkYrv3PtHI2oj4t7laWoYl+1tIMgPXB+NLS9NniBwIR34b58nESI1vxd8Yhhm
2juzuaXoJqFhfWpMS8wgRcBn00dKpcsKyE0b+OuSmM1JOQ81+vGroNEWpNEAZNWbBqYp1xKSXKUY
/We0J+/PrgZWvjhzWMwRwxq3EqQ6BXjHNtn+rh5RLS+jX2ujYhg2Pvq08HNSuEU4jlKKlEJKwfL7
fmj4vi2rJjxBJ7eKvVJWtIqn9CkpcjpECaKHukaF/84TETt+zudln0T5/90RPVqLO6crLielyNpv
TlPD+zJH/shYxv9dFTWOu7uBBKOdK767fIyU19S89Qjs1XwZzF48umUEiwiupEq2tO2O3/yxMyVn
yRJG7DAGKcgsCZqOiqQ4cmBUQCKFs2j2FtmLofiK/6CIUODt74bwtMJvaA53Jn0bcw0+0uHkUnFt
XnRk5qw3om8hk3ZLPLAT0q8fEfEE1uY5W/eqz67yuqODXY4hxbHKqj+YdaPsoAWPczADVmTorbJx
s930cnk6Sgczd06mYxbLH8qwHPPxef5pahJKgxZhyiTf/ILmWGmHLznbwOfKYOy7ki1XiGaRqvvr
3M48YPHsWaYtU5EKqRCkUA/3lsTPmSnVku1LVaw0NKw5W4cz/uFU8R6qtDvODPqW2qkGxZoTncGS
yp6CVBnjEds1eD/NtYEwDHm4X1LEGOwX2Jb052JeTbO28HvktIQiC0faibGxeqRks/1zvQHn+zRn
01qGIE/9N1Cx1tf13OxanwqZn0GLbYr/GjTIlP8iLD93AMEJbUo5LxzHBSNuMXOX2yLCO8a8m8R1
Ye8STwcvv/KFpUcslO4pDnaIZx8WT79dnqUPAHzi5EUXGDaEn/cs+/nNNd1/NfdYibv0lLJZDHUW
XXMd7IPN4E8Lx2KJqpceuXPiqsADBhIRlTWnwMlzwfgW/gC7AmBjq4PgBYHmagO1GVU8DOK4zcDp
J2Dzb6U0smzLxYY8f1bx7/dokrpuekjrhhkVhJgU0HRlp3s+UlL10xPKt3cR3KfXJx7tkPdx9vs+
2J0otF+0ih3R4wsrTfHSCfu6Ce0IC00gViiYkmTlR/+IpN+WPoQ7hQdnNeKRwCd/zxMQbjghfHPA
agfpEqrvW6+PMPBFI/vD5PcXSbQ324d65Xe4Stx+yBx+oOCkL4maMYq0aZQQg571J7gKJQ9lxnwU
TMH9xP2VF0cyLkfmTl+JWypVjE8J36FcfGGw5fVfGPb1ric7sfrjNDZq+NynGD8jWveGRFNYYYPv
TSsdSrJnME6pGUNuAI2nv2DMChEhhRNw4682VnjSAlqAqXZZpOqdw36F5qopIapVA0TCszxa9vgV
gTc0OEJrL6RPlnDK/HBb+fO8beGLBI6AALu89GbAb6ObtFT/JYhFqiIsXLOjRh8VSSjUItznKpKS
kp0dkWB9ozrCgmhfr4MyQ25Nsm8/TPWmfwbleFgyJFcVlR4+OatCwOS/l2AeKfG5MwJUtELNDglW
QFine7ogVjsQ4tyA4TI3iqY7VXA61gQUHlS+Ld5TpeN1/0VkxsJVpHZJ0mLKtV9StJT26ggG2z/Q
gfoSqu2SWNfVrv34cote2hHGbacRIWFKNG5x9f0XW+zsTBD+54YY8K1lVc58gUeJN6pfelo5wOq8
LFHvt6zlj89cmWFhG3UiUWzxg1BiszMC6I965MsxQ703SK83N+nQELwqz5xTK+HHI5Pvch+O4SVv
Szititd7sDzXoBqnQogqHE5Rvr+4Uz/xBwFFJDl6wKwkbYF3rWRLW9WBD8xdUlHj/fgfjzqGWNe0
h+gLdn/21oPoI3hPFU5/qQ9D35yzBH/rlIbw4JPjl95KNRb4XTmvxpQo1D3Y81Zl2ibdSuRI4esW
H2sDoFqOHZ6ugw5Xj/Abuqn0xAxzpikAz50FfHaTB5C1uBowGu7dgq4V9AMfBG5SUhJgXgTAPYXx
B2PZ/gqpSwVMBmaK57fghFOnCfz4o/ObgW4XB69QKtAXz2VPPQh3EXN/bQhp1txI2g1s8RwP/aEe
PYS+JSTm+JVds4xFKtGpsHLHFm6vLMPySfLru8/azdMGeHtgz3OXgb5qJSrhqOajmo47zbvSw3M/
sO93trPRDUpxYTeBnbhx3hdBov36x6AExoJTvsyRg6vKZ76iakLS7uk/aOZs7TlKLQTJNpr6UND3
gx1oghZH9DC8tOD5zwPQLAzkEpyN+Wb5Ric4GatqHbwJZ/QDwo55oG20ZQf7lPpPQ82f8pqau6Zw
boInUZQgZ1FFejY6zWymvb5shRpF2IqE+VENuNHr8fq+751Otn4nc/oOyq2P+gH2RHvlgKZMHCo7
3qVYFoaOCUwD7YJu46bJtrYLYcGFe8S3srJzo9GH9tvDMS/OlAgjEOezJsDyWePU7uJcBmVQ06k4
fDGBtr+hlEGolGrfHfGVUnJud3L1dgX2ut4EibRyWJp/4bwf0xipmJUEYaBZSW8jklkxnc2lgkRn
d+BmcSRK7jT7fo30tdcw5tbxoL5SStUc/HGiKajtm4nS6WsPVQvywXeGgOvU2eLfjrUzJ6vKWYyo
pU7eWGbNiY72CBuCxVBgwtV8Afe+nX0839pnPvf3MIQnVA82l2ZA0FxD7JXodacMPssp6rYLSlSe
QYdJmTECTq1rjToS+NC5XHLYDzvskFZ12pbjPUEoFhXFJBMbnDHGDMb2JlU66MoX5Z/DFUtbZJZC
ZKLc70qEwcB3ARvtY2VULBKMEoa5YxYcDA9lVsiqRVn6WsnRdekbkvXozEvu4VQYAo9jVWUbdg4X
a9VxDiavd4bkwbYyESs8hZoGdBy4Amg0M49+Rkq1R1lhcLwR6TTz1E+JDeaz/cPL4r7fbPgCn1ID
gt4PgaqJnWAhT8ds/pKlF1z/x7N/+AJWaxYrwm9SHRa/lIBdoGdf5fKm3ysVbQkjYDbZsgUJthba
CD6weCTnDPDMMJetu/F9nnpxQmAL6WVavThyZY7aGcN8fvXQfSL1sZJkK4vvWUHPgMd8Ua6irShU
6zz1dc/xN1KYst4Ri7WkOSvWTYRg0Gc6yRs19JiA3y5Fc7mNgQHLqR4Y7os4+yW/WhmOEuZXqCIj
ICBRlNjnvjM7koQkM4AqtvBLDZ9CLK7L+Y1xn0BGrXdHXlwVFYAMJiBOSwuJMd26vUj/cVRHWrSQ
I5NYwHaAiiF9zKHjK8viRmDMDQ3EY6ebctOx7m//ZeU9soO5F/lp18Ewtpy6qkRzx2qsVcgXLTuo
8APKALM8zfmcEO0uHJoAkcXnOlv3Y7toOpDOK7nhrAPDSEH5ZwVLgxHcS/t6EjyH+TeaW14y46CJ
s7Yq28B4Sq/zJwCpR5zUKNlDJxJqY2UMqRktT9+/qLGN2csNSjrloSwNdH80P9PUdfUovoUzwucJ
CvBqim5cQUxBYcp+5xtd1FvN4q/RKE7yvuNqMqKDeBMFD0khae1p+AOAwIh/a4zZUhNyEvQgMIu4
AOCNZ68kEKg3bM7qkmvTwYd8B6ngBpfnJxwmnxSSen3eM61v2zoei6wgLSdw/fV9FyzdKxrlXdfY
WBzBChezZEq4/2q8bWNVK7L6f2HLf4hum3rbDX6Qk3qAxyFNUP/3yc9NyNwUwY7YSiQJS0qbIwR7
wq2SWL1DY+d2yf9GOmhGGCz7K+OygD6mcR92tdj6WaByoMubecUSJzhna79VXbd2TTmkhYgeZyA4
N++ayieLpXX9U7zF5sHSXuv/ihetR2dKGlWTCeGhAlk6OBaXQDq5Pb4ASEGWQVJH+4X0mt562Q4p
LBRommpVSM/ptbwQDwR2D2jviaygVru+wUDLQV1JLeKBBaVtiC5EGozedxOXYCAejbPm3wx+vhFd
3HpCzDz167KR/zdrMSDtIV3c37z1i1MGSiJl19sya+Y80ZWBfvdNqD0sdPY7BbdNIfN4fEoJaWmr
NTupILqOBiVWhpesPZBHj0mvQqOkG5iD/OhkYd80idIGt7mmmvzrvdsZYfkqT0wEPCAgv584M8q3
6E8VCLmOyqe15z11bgnYwOql5r0GoNlf4yGYYjrK3bUae78Ko17uYgVi8GHYpOymaGddSDOd+5vu
l1Kk6DP6D93jrzbHZGNxLz9gGSI3mzWAFvJU3bXFAT+2Oys32Vmpbgpx+Gz0ywoTWlE8nqq06c/e
laBEVs+HwqhWrUmBewmExDFw4NSJq9N713FKKvfa8bINH2GILL4D9Ajr4RvM90354RI4Yhoy2+e4
WxdPwsyPdlSy52tfjEJEoN1xYY7YxWMGuADnlGEEGzRJ+iCvv9IeLI6Co5ewy05tFz/+mUAKYYEt
Jv56WTjDSqdgbNiu/MdkQSWxbKK3S6R9js2QYGLXYIvxcVQRLp5NT/bZrC6d7VTEuLsOaXzOMl6F
h0oKn1LYxYIuHo8TXBFkJEZdT2RcZETHz+Fs9aumKExRoMJwx8YQmcvkhsHQlR8bNfdhe3c8/ULS
X7+95giqdaRvK+v4yP4a31pqGXsWKwuiONOkWFJrofxkJfTp5sooHQLTih4KzpGr3Ht9nyn58vAT
PHuEMHD1rWMMzwptiuz0p3yuYgsmZh8lJwr/EhEdeepXp8HpcXoOEEkLuaqX83Vr/r0s1AE5zOcz
cCBPRZahrc70bIb64b0EfosEOOYkhlqmTaXPqn2ixpwxQ/aNzeRKqkZvLz/vI6jkw6MBa+uZogzM
L/RSFpek1+7JixArtgA5ZRuHJlP3ppnlv8hFPMkUS8AG8dHybddPH7odnShUNzVylfzGweeDKAX4
VKkvrTrFbLRQKmCtrj56nACeT85YohM11oM3HNSNTfkAJonzDWpHF2yszr0BEn9eBfuHzopMsJYW
a9f2ImV15UEgrCzOEggpRaAgNbcFwEYmM8/GJ/4+UeWjpB73SYjETR6pIE0YOz8h55RJpP4cbhfb
J7iM/rga/aj7ps/uP9oJgtm0EWnybPUTV44L+C2/GQ2Z9ZIXMrYk5lKyw4CK0j1JxNSpKP9ci2vj
/ikZzgjlZK1Jyx4LVOlGMgIIps8KX+CrsqjUAoEuGaRL49E7s6F3HCBASLWz/AWsGFJY2kUqw90l
DLowiuGuiI4+byENeoG+Psbad7R8eONlWyMFXDFX7S2x19VKQP2o0HgRxgm1kKnz9G+tBd8/lgh3
2KUxY+tze0DkEIq8AOT5C0VIadLP7lY6Eh6Q05JQ7nw1mCfEIhbpAtEk05l/n2SQAGlkjCxszUB8
mq121AdmH7XzAmme8tw5O5PXF+YGmHw5S8vzJNKT2iLElyjv1idiXvxxY5yh9aAEpnTPfhsLTkvh
A2YEnRUZtoc5eftuBtzdANfrZKImj/Kq1E65nYv2n0R5Vhd+HUfJAtd8cKn10bXmPjcSOwq2So82
cKqYoHA01NjfQJpSNiW4iMb3aLgpe7lVpgjpKFJumo1c5Tml39//lhYkRoRUUYNrtyPJ+0TvRQap
n/hFGUDwySMc7WjNNqLm9/b6LaHZTyfWs5Uy/BHgIVEWR9p5Xy+78jc9adaz536OYldtv9gYIkhb
X7jWeNlIrJkAkSlWVYffxe+mgJsGPeBVz8mAeouVfblqUNwvasIKut7MSb4oEoW0W6D3wQkKlteZ
tNvy2mKsun8ykVaSRtSZmPgkkYYcXNhcegSYE5UMSshmauWO6Krf7xksCCBoFUJQI0HG4bY30ycL
hsezPna98kU8ZmfODGQJq2fWXvfAnr2wu53cc1kaurhmM0+Y2OcZpBUKbHl/bGtDrZ9T0FCDW2wF
rDkqZEFTU0kL47YtZ7UF87GjLyAYmBZuHztJATeHyNr3QaVre0aGPyp/TDL+CT+IXX2e8HYG0Im3
P03JN3BhRB0psGrkQuVVBmWbFbjeNSKTPjraSORFh/ZHKgyPhuG1ro8+0CxhVqHbHTitLJNRQ2YF
ooviDKeztbjFCtYacIRCbU+zsqa2aMApkKPSw86lDUv4rDp3jnXvKGnDe/O98tA4TeJqVtygs68J
xNYhUMkBzhLGcAjNkEqrsMgCCC4914HxSjVKNKcw6Mas41/62b+3I65K1449Ah4dSaBmLALNRcBj
pUJVEFx9OrCJXui+3UYXVaPhiWhnMS30kpXFN8DznveY1HImTkZVV84HQF4wrl9uqmIY1WhoDXD8
W03H4NoWUDhrbn5y/3/+IE61p/c7RgkFuvwKPQpSQhdBCnex8amsxw0SdV3Ga+ctQsWuelcGT9BA
EBopZsYaizWtnX10Hly1JsX0zJ4qXacDmPAdFUjpFZwh4Q0iqXYBYBiD/r4q5Ps6TryR4+VPCDFW
/ulKf+hYSZiEwj54e/Prvk+r85jS9I73a0ANl4RpY0Cukt9vmoBg3+G/4Fz/B1bB2WMX6dXg+LL3
sUgTAT5XVKUIJzk512+cibT0Au9xlLZcoyKkABaRuYr8qrobcbp+XCA1iJl464wGkeeHFzZMlpwI
6WF/6cG+2zpRzI8TnWUX0U6C6flsrInl9gCmB3RkA3mFdWc984Dj0Y9dHFh+3MrTnepCktgFu/n+
OckT/yvFFIsiKXTAo1DZndWTH/G3FHUCn0P78fNM86vvbEYSvHZpbPWBkzEZ4P22gJ00yzZVw3cD
nv7DOInR9eN+ULncUbFqyzCIaYaneMs0kum7uBCSj0FNGbmDa5KRCkq9t+r+tzNsp+8sQ3od5QYw
KBiG2aK5th3z8RwQ5taeU7WJEkQzU2BbrqlvXz8bOzXbosRvgOPm+go9/hr/8COoprSgiTL51fQQ
YY8kWzYLwdzaKgqh+PqTY+aOqijnvQRUufzi8QZC1c45a804VQOkItb6v6h2MedSS8q6AyD6H3/r
/SUIFy2BB9oUQJcoDDOeoqZvOdPFI+T1ZHp3cRb3u8s/pqFB2XlI9182Ix0GwQJu/g6wCwSaAA+p
+SgASsNO8yDa2Ev0bqX3uHKkDU2vPaT/bp2y/MTUiU27UbLIRrkfRlpsk1wpMdmQzUkFwKGesW0+
D7UdkHVUu1Hf0BUiKcPSPKDxMdBzCXjaxdn/SaqnbAG3qVBk0FwBu4mhYZ92OMfW7qkvjfiDKPYg
8gb0KeSjh6x0GbvItss3IUiyC8mc0ekWtpBG+zMl74kRQjNRpbPqXmvq78S2v7quzhGgFzUedYL1
OcqJBUdJxC8JSJ93B1Yllox8vYQh2Mruczvk9e1s+blDVxDKKhrmpg9/taJo/QMRuhOTdzHD/vzW
dkNRdTi12MZtcT5QLf4I5UnWtv2Jvg65j/oaMaX/hl36qGlfiltwFcgcYs5lITHOuDPWdsKQCuc/
P9r4v7+KvvoeaMaCVCtxwZ4WV9/RZtLkcyrTAnq4o3oi7bMtxEHpqTXaTiTH6d7P38YA7zc0o9Ig
3AGRDIUSqsAg8D3h/v98t+Uf/ZcqYTFQPdGdDEWgDlUfzWy1KJB93XB3JGiK790uLq6Wi484PDsh
y02d3/cKmKSQRupRUbVVSy/xHGa2twC+wS2e983RD8apMhE/5OvHlGvOT9/WJFgHdaosZgvRvbNL
WR0qjW+XnA3TdKLoFmSNR+pSlSoYmCrhISrxzWZF3AZA9iBBy8we4Na+zN0qHlmEAUMGzsD6gZ2R
kzYo87W6YHhFRDIcDtj/pE8RhrcJrC/3zgvCvkbDPi/I59elMz8WOe7QusiPm9GVEEqH3vWxq0Xp
nY0u07YRrserGEyP06MKBi5bMf441Drs/ZwCpHslNW2JAd8hCuV0hjMCBcPyyhEp8+4HgWRzzIkV
3nAhwRod3Z3lrfM8l2q2e57mzAJfoRmbzqz6bxpB0kz0kaoXoAGqh1LNVa3wJvtDeJkTiPSeiHZJ
Wz9ZCLA1zcB7nfVRj6hcjwDiQdF5lnLoOmrf7SmQTGRsmbnagDtgKG5kl4kR5hOdGBhi5LmuygeW
j5E4z0v9cxrjgp/p+Lfe0R+MTKBJRfG6V8DDhuPsasale7ef3y7DyeY+lWg8A2td/imlHhSkRCCH
Ki190oLQnF5NgEltHT6yL8RV0FOsVRXhvh5dFtdN5Poy7Fbe6J4/Vuxo1ULtCBNip6qTIfLWwryh
kIUoWKz5RPuK07R9sYRyE2Cyq2/Y47saDHspOA79T+PT5SxjF17V6MGqET/ZXTSB8h0VWqbo+dWJ
9FGzUUGl/ukCh3O1iiSHoR+X3mFVx3B2ohuLZ9OGPOOlG+MPSYIssCazAru9x7FTW/TJyg+dBUzH
xAVnZ8XcOcnAiikZzUt3UfWYtpUsA88WnIWYA+Gm0WZDpMDZQVg6xUxUu/PPCqJp/aW/GwlIQTUS
nclD7YZYi13rMquXaw/ppbsRbgM1R4SQA07X40xJ8EEHFNc9iHpLi5DhgH3Gwgt9dG2GXY3y9hBW
gdnJYWA0gInMYWxujZ4pvDonIO6VwRGGSX+Zz+euO3P8lwxjcxqP460mWNUCVNpFULS7kPSfG+XR
VOWRPKpKpC08Zqlu+QSl61wNPo89PhRLxfTeWu2YQMrYvAto6L4WW84gKU/ZRvV+oqghqDMzQCmr
yRI03ptdOC9NtunMFV1729tvCwkJyQT/IGazMklCfUde1NzO8DspD6tcPDy76viomX+U3XCBaFVn
6l13rKisw+JnKH8F3SQbTleV6QSba3JEvAwrAV5jWofSmdzx28x5RKrb1ajn/1P6P/aLs6Hc+CKQ
n6z3ypB45XqS2LE/VqEHNAC5ZQXkMYtAaIrtH05pE6+yqu6d8WDhSDVvEMppe1wjR+b6zk2N4ABr
OhQNAfYE45xDNQqyurk72RH102XjbixKK2v3MDuDxG0BlDFyICPLcMwCN9W9O97BeH5Yx4AeWptP
y7u2haQ+4HTxfpVIRJ5GK2odvy4V6jL9gK9caGiWbwTYyx0GDAmMNYCcQ6TBRR4W5foOw4CbmexZ
PMwuzu6ojGBIq1AuJn9zG841n6Rkt6dUmrDPrHCUOt/WTG4C7TYKVut7XfPR+Oh9owdztm3EKJeJ
aPDo3IGBS6Wl1jiqouHdc+QadtejLMJd1TtO2MsldJemZi91FPH/yS1PqisamTs3AHW6eoy6Nj49
0Pm+e09NmzHpOGQZluNbFTS4T9g6guK9z4JdG4ajJBYeh/xyJXJecLxQJQE7v6IbUh3LzKFKVbeg
zg0EVoo1nhEOSglgrrmhnvsJtZG0r9owBhjIAlfCNj65Ub5NHYkX0s6h4jjSuNmzgR/zuvWaEnhA
IMZD57wP/VR3Y0S/Bin/lcEDrtjIOC34PHQhamklOm/FSY5I/qRsCe+b8HOxnyHUklQzKFZsb6CE
9JQ6hYz6cMitG1Bie79JrJHqfYeCGpcwFfaKB6hcuwI5e/iDiUVcIiBAP1tq/z5yHNuk8c3QC2no
aHeVNrsbtG1MKxHw/mCRT82p+ITlRgUkzHwbV8yyiyk47wSVG3qLTFqfxZOavNPHdQGXD7Kpk57H
um9uQlc3fb4+3Oy+YKzJK+amfv1ES8ufTkDR5GagZ2S/hG39YIa828QczdZSm3bIGnT34O/Q+HLu
hoHTi4vV5pWvlwd7veSd9tfDER5uqer1J3RDiUhgZJ1Z8JN0EXE9F72eGbk77nN+9UtvobnDuXb+
PpcrkKl7aWwG242hs3j6SEiLwT8q4dzO8Ww4hK6e8qGiA9M2HDy9MMj9yOC/L33UXMz/MfdR8lYi
vncCTnynvwdpizBQWaAZ/tECi7/J5RBCzUWPEb+CJmUz5tAER4Mzqo491ESetYV04+3vqhu7LJGX
j+UC+qFLv0f3wSzb5ZcJ/SnVbCV+o2AlIEQDIdy5bcLIqOIF3NnigcLAd+cd6k6r0+riohrtNC7c
5BINZFnkN8z7caLSfznqLnJbEQSe5qr9clIVAs37ZaUYBc3LyCsqW9DgAucQBxwi0oa6dKDyulfu
ZfdqE6dS4WVAK1kXHJ2qMYYS6jhsuxVTX92Dap0f34m6x4U5kk6aL4E1w/YMdGX6xedAIfLKtl9b
BNwAYaaIVLesISA6LCuEScJM/d4BDdoARntmmWaVGv5dbhkAq9VnBKsJ4I9ev0lwkdUVMu7OAc7J
z+852Iw3W7+9d48uO+6JflBbKm3tAy44G+7UreovJjyGL4AmF42VUfIGdI8/Bkoe2AyAc7JVY0bV
bBXHkcYDp5RQijeVda43sm8ylTzeodCcTk7ygqvZM/XOWFZMHvKVIL6ipU0NZZNMIAi1ZkaN4LXx
CMwMwq5yVlD4bH/PCnFMJ63w8mzHztQC5+s1cvi4lOWxl4yRBKFisNP8/YyGLIqYcbRl5eR+Yp01
eh2lPVMyoSE2VLzTM1mhovgz5TWJWxfMaXe7plN/t0D+/CYSayVMFKcvRw40+onz3zQLOoPHrQcN
CZfa9NyatBID4lUepbK5r6g3Fa0LFwYgmkoF+zOS1+We2+qyHiPSFXoZ4GAzEUvgxZZlVDRJF86h
9yE6HDEfbpoWg/Uvfb5NAsoCeyKvpY797arnBSsLYvtHof4FNnUuj2/gEI8OORVI+5DYp0UdfDic
a7hMICo97oLfmIISZlD+Ae7lqoQ2J3Gjph4Zn2HJGuZvTFR/ezXmR4tmkz36QP8sorNNVyD5JAwc
YSbNfqa0w+xdS/vr9T9hNqqTiSUnrf8WTIUQyeAq/IO8sI8aSZIP9vbaXWVAWLQsPmcf1Jl/8lk0
tXjub/sT4rdDzmcBkI/GfeH/d8GVvcMoBudiT9sbn2CwCec4RQ5tVNUsgvmZQ5Jl0FBqCuwnGXKS
dYe4rGZEnVx3/dIps9KJJvHwyyKC3jYHlU7mdJJaVrG6teok2JmSvTDDaVjiHBNZ8B7NqpPXGmWQ
inp1tJDJPufBglp3+E7D3XKi4SQlX8ZjJ5HM30L6u/Dy8CknpCjskC87ldU/V86KkzaVedLhAxFS
4nI71SFZT8Zj5+Qbc/oaEZWcwDgDQ0JXXml5cScw6oGwItLRn5wJW+szYikzNzLbioAhA39FoP8M
wT93NWYwsZEpURGLHQKs/k//Pg2K+gzmgF0fT77pFuwF+1PlpCk1xji9DxIVOB3GJOPPQLSmU++U
QH6jtEnKa8+0ygDudCxllWQt6yDMOzqjOn9wcaTH+PO94YkRGMWzgASF5uZucA60xCvVpVLl+m0S
tjYuvT6I14A7/rCj3RaTzb4NaIf5Fr+zPVhrRpx9XOt0dH6yiu32jAjHDUhuYW8zi6kgXE3Trnqq
l/1I5/ia+UFOQLtAGXvDI+l1fi1Gs2Nx0cFYy62bppTm5mqYIX7Er1zUWllf1IHvYv0MCzunD/xD
i3/0PRp0RQVmFQbjVklT0p+Uf37sTiZoSQAJ3dc8xCP5SD9Ju0bLJHob2zv9Yd9BRaUmU2p8JcGz
7DJPWGQuNjBQV9hWviNrx9Mf57njZoBxFerHYJRFp82U1oMNwfHGs8tEKXlVn85AD3yCdEuDfqO/
Rb2rV/xMD/Pcwg8cULp/yIkG3Son4btiZ8aMEKEi7vkp+a3XJusQt1SF7kGQFZG0YOP++6ajorje
I2SUiUCUQEwZeTMn9+WFb4vOcu+opD3rVIWR76BcpUlNaZKMVuQec5P54cFvBACaC7GvJmwQcTf5
s5SFcxYG+E/Inbpvj7mKPIph7K1D5qmQjFR34Wm2ppXPOahCpBOoDwBCJZqcc6XoBapYFuxqmM6C
q/E0eBiRJDSLVeWVEHrLFdl7ubims2lLqk+KqPThEfvhjnWMKV72eiK5fdE1NsV99a3DttjxDY8L
L6aeuMAVPIZ9Ry+L4o6wBy4NjQa12ekZVTcFPNIL1HiyXOJvCn11N5GndDfwr72scM015lYLamDs
YjbhJRAELifgE3eZNtuuOR7wKz73xOBpmWHCqwdFgd0dta5visnxCPlz/O1yzE3jtc5EcVq0qPsg
kIwIH3qZauFZPOnjjxyTNIQViOb0ps5zROb6DNcnu0n/7uejrCBjya+Xvdofhz68oVGkLErrw2sD
2pT0s86aoQka6BP4GkMgkiDYyvsPhgodR0tcck4M2KQNUqw3cn6mkycTaGixiQSXsPVVQdsw5B9U
2/jO2F9zdtTYiAY7udBbBfgL4EcB2j2lNCqe9GAnFAJnz2M7nb13KJ2AE3WARwooRdVYEj0brieB
perY1Fo/GljqlOKX3f7+5PDWGWTiwC+Ib67zNfModmcNOBLh7ch+VbGBQMRB0pgkOMpTlJ2nJDyX
hicEeV1lzGplvd1K1crHudq5kXIb83abRm1hoA1CVlmEu071R26gEOMs2JQxcysWdcGmmu/3Lr1J
az+ReJbInRzs9XPE+Bw+Tmn7dum7EblJLTV+8c0lOJKcGmk3ntTUhXRlVcH1NOdZDJNs9mv6ILTy
wwdtwKEHDkoUFS7+wGbxmUjkarPCTKdvW2Q9yjsWCmb8wdpTDwt4GTbuHQzg3C8t8B0WLT5yQIOa
9xo99U246kWA3uO0fiMHuwtPy0QZCjWBWEEFb2hD3uqga6Dy0OKp1KHLs4XOCy9Zrv3cZcA3Jnub
bQYBrQYJDG3lvcDJpp3LIUlDtP0zS1ZmnPntnIrEL5Vx6THJ2V9mWBC/y74zYZva83gQOKQuSpAG
azNBqHphquaanJnL/De/W98Q3y0a1I0F8ZHDgkrbTGSASKeeH5s/5d11hy+khb/MCKLjEimFphME
0IrKx6twOn+eZ3IFZYo1Tw5MfGMxUCQHCq5cONfqOuMWndCgRijGS2HCGWoOgTZFh84DPm4rO7VF
m2PYnYNx2wXVA9SehA5ZImXr66wg67S8hOOcWKm36S3103DBnRU2CsPXVyFqax3J0DeLupmiVD9A
bSdt57/5zDvB+Qqiphg/dK0HKpx0PDkcTl0ZJerR8OkwcU6p4D6Zuozo/K3hiovPCilpqRlsepEm
/sAz6lEN8s+WhumGze5jCcrj2O7G20u+4XLPoiCc4sAivsey5rx+zlQkBpXV8Wp5p/c0uvjaXcIN
lZtl03f3BQvYjl68l0GSnR3NkU99jXQPFjKBN8/30RjilyeNX9/RRqadOxEEJ5YpfqUHYztrfCcH
LJRHSAKhXyTrst7S7iICjw3rBTE+Bl9pHSAIkmZ7aTJvMbVHnwwesd1qRSyUqZMpT6hUrGDmyjkU
q1zDsKORM3VHuYLEVEHOKVuLLnmqQCHFowH7CYhqAqDQjucGm1QEcVLuQhME8T7pUbTUvJtNWMkw
nIy3iGnxK4knEqbLDbs4XkprIRYxMarCl+JbPE0EsBo6az7HFrl9iplxM6legvLjQwqFQjH7omVF
UdP9VLGYXkx4eXtDplY0rjeAdZ+QCSCDV2sQDlvicjdLkCH6Mfx+aFGY9dSdWPzqzODtnr3kfWwd
izSysWH18tp1P3L7QKQApPhEEn1mmsclGtBdCUErXzAMzUHw2MWhKY48Nhknji9o2RZ4hH82ROBr
SPv3sB5gJAjami3BdrxfZ5s+Q5ub9H9S5lv6Hl5SvYNfcK1fYBqe721oUkDIeLvwd5P0WBgmF/g8
TM39TMyEwQbnTWXWKkaQpUpdbYnID/ba3YvZ+zvUAyQwXY2bGQCvpJKRdPRL4qo+nHIPYIygfpSC
dqEQwIiGNxL8LY3AFnKgtoSob+JaEOwmUhDe5Qhag5a0RleSPLprs4tC8skABrblMviB9u9mOPfT
XVqwk0lueC432kk5QCvcNyazJTchACGueP/agqG2CR3Mh8veiNCdh8ODMZZxfRRDNALV2wnm0THJ
O+VZor23rMd28xSMXAjqg9uiT4WM8+3a5o8tAbumAl51BAAlW3iYr6+BqpT0CzmnplTKMMyC7GGS
6nNSqY9qASI6X6nKMdTqfGOdA4y2RRM3wlLC64CHYarcHkHEYGOYbZgneD8Khp+81eiSqYZIfAI5
qkrrwgOswUA6amm00DAKCaH9WMRwJcDh+Xsg2viIZfAH8IaFez9CWRrahiA6lWA/7BZ8zwtIj72Y
TC7YXpiHeR0KmLb/owYg5dfsLKeazGLuXYlM6Ozws4mWP+FhNZqVCIgAXP2rGvIy9UzTq4L3K/Qc
FJF30qFNAoPlNyPivHYNCY0x7u4ALZgd4LA/IKo2ojdQ2TNcYMvPKCLuuohtJ5D1JuTzk+LwRvMa
SLWjFeARsaq1AjwP/eIKrNHXermXl0AvLDuqKQermxwDp3s6A6nf350TFAcnKrH2Jx6QS6yKecn5
aqVdCKdmhL2Q730a3+3XS/CUIwqMfGsfbh/MAFWtBwLSYSJtHu2PhYWMD5Cu7Kxx3pIc2EXOUm05
R5MvnbX8LmGTrFOI8XOxRQS31lBcGo4ROk3xPM/zayNKChozaKNDknbF3Pe8JbZ5ilaL/gBow/cQ
tpOq9UVE7Z2UGFzrRCV4qEfP6yjef10hr9ovTNXos6qj/YKh6VsRWeZzUYpLwf74Che/IeHMMMnA
zyjkOzxmpn6yIxheIwiGUDjz6G1crB9K0TJ5dOzxOUQ35Q1qLrd+Ejl+2m8tP8KJdwDvTjMby6XE
zLa+CZQBHqQB92uMXOA/UyRajGBe79rQ5D72FUvgBqp3CFxmPoFcmZ0LPoielNPT8vGQ0o9brZUh
+NPEKBA7jRI6yw8jffSpBGdL1CvkwXrpzp5BHIUVoPgvaTmLEFR6lMdeM1tri+EyKwLpvqG2vYbl
78iSn7SWhM2GCbkZpn0KNjvlXche07bXe+ImyOcd9Ep4UjLFBoO09/JVTu4Rv+6KuWwsFon5RlDX
fS0jFuwABkcwCwPvQj7ew8vmJbcxqzunSTSm4fkn3n9bupeEY1Jc0X22cXpPkMEuCQWSELhlyMt4
mK2a6uf5u1j867V5bR1odvc7Yk9giT7yVGYampUsCY8KkK+iiO376gxoVRtued53xeHPtRTNU/jI
Q7kn4fPHII4+VwuahqFWZmSsPwoaD1rMcD2uW0VKqFZBuw4nN0LSa3B86W/Rc+HKWpdgO6izWPLO
3hIsjsNAQG7oQwpI1mNCGqexj48Ue2bNePV9F5CDtF/t1Ofz2izS5wgfjDV7VcximPHhPcr8aLs8
voFDpAOjdp0wfkrt4t3KHmZhF5Ju1AqD291Pptzf+QIVXLlncsihHpiZtBbM8NMhlfQYh915fXZj
PZLAD83jauRmqZdRObhiQOLngJ0fivvQt/Jha3nt8VL8o6Mmtev+R9YHk45q0qQVEBhyHKCglWMG
PMJF0c5z+oVU61dK34VmbRsiC2ukQ+bpMNv94CNisJPUFfY5hQ1yU8aGiV9avRHBAM7DzkdoqEEq
LOkZLuVIjZFdOl5gko352ukndsQaJm6tSHO6ErDpS0n8QRl31nf13uQQVpzYWG6GWrQ1ozBDv5G0
aMpgWtO+FohpQbrA37RYwemsnSrX0iH9WeKAKd4/JTuOk5KN9fWdsKGqmWaTfFweOK7iWmTioLxk
GtKaWwfdCVcLqzyqdrKBDoL28DQh2qwvpxLnixcfY6BQWzWEEUSj91NzX5l5Dj8xjAwPmQ8EdID+
C7LBFDjjDY0qyzulOAnxLdZYDFbWReU/+WIccj/9XzzU+YNdgKGrktMpEAEacmnAJbyCbgLgtMFR
+Bag0ANQ/i5fQlGRcNhh/thYdVLdDYXEtP1MlBePZIX0sGd+INI63nw05JlHxmNIskWL0JSHJ3LH
2g/KbThOuwGrumWzOvvntzXBAbtMsfs4v5UspnQ3P9i7CGvddNoRKb3txUMkvUva46a7nq2nLfMw
VsGxYIdxSpsydaalLS0VojJhgZqDdyzhp5d2zygZL7hjmi3QXarywQT2BN6imk9jDY1c8fteQ4U8
ATVRjk3/VPxvNZYCMo4XI+gjhi1hCdoDvSijHn1QkVM+sUqwe9BHKdl0foxoHfkPG1HXjYVFoO2h
W3n88Y+RRmzgqndYWAv246Gp9d//zVrn9LoM5XmeqBTFwsky9yqzm5C9+qOK5gKZvKpim2Wi65zC
Z523oLE037dKKfJhF7dXObBYHpT54ACMa4S7Zu4JZd9YxI5pmKWxy7FvjUrINeks9QD7KBKa4Bs+
+5FDBr5X0m3dSxBIqX4fpfsyNxro7DWV80dDZFcAu5Im7Obp9XLkXiRbidZ5tKJxaAMFN/QF6M1w
KFYX2rr6ObRhpXJ0n3aVhBJvf/S2aldcBF/LaEYfAaxEzmV4uMlqegW9JRo/6mZzPCi3bor9FYPY
RP+bS5JkD9fv/w8FCNnDU7uQCt/ao1jd5Utuus0TNJ6UHIoZzG1737ntrhxXTNWBaEOA9XG5WM0h
ZejYE7UN6QYkvi1NGqkVXYuZA2ESvbvkYZtV1+NYVXuZPTTo8/Ol9fA7m6SeIu8a/v4kqQL3rFMG
G9sHfYy/tSwjJnlNjwexjjrCjVCadPw5xnLh0iLsdzPUxoc3aFAUONFzKOQE+x4eLa2H5heHnAay
TMRPuzjTov9wPIlpOSP+BJt32PlPWcNW+eTQwaTObsVq4Ix/V5+H86boI9D8NlB8GCirhAT1tKKL
laHGchNb2j85rct7fjlCcWmsYdQpKWmV3UThgqhBqN8t0HP2YXHcKVKFtNfC+xfybyxqaUwGyPLx
V1RElScXLlajlfXJqZXZutgo+82s5qbiD32UGTyPaUCmw69Al/oJTJHCCNdB7XZGzW9k/7k/MYmq
D52eQXgqfk3VHHiDZEoPijcMgFGzRhwCWigPmbnoExdW7JnWbq7mtZnNxXB8biEz/dumhyXmur7r
k1iwrQN/pFQ/wU7sY/26s1zNX4ItyGUtdoR1kV6HEsbjP38liqJY3xEPLqSuA9OKQTnXs+/qlPV/
Z0VenlPV9HVuib6G0DDaLmHqznJ1sQnGuoMBe2tna7cHh0T8/oEXbfOq7gmQkjhjO7EawPvgn9xB
n/wHgLl7kK9nRJ+6Pnw0ZVJLVL6tDeI34fcJkNnzs2bFksKoB2lvZMAr9pcYM4yvBZmA0InoI9p7
Fc2f+60rSP4u/hvKNyanLHofq3gRJg2X54TcEqcxjJqfpqHqZV+ZJwwSFX/A2biFv3GWqAkDyxqE
VTwbSgqCYCPEmn4g76pDP0FNlDSEngRR1Zs4WVBtytyaGgMN88U8b4EWZ7eA5Xw3n3K+Iqz5G3Qj
LdJ4s0KwOJptEAYYe+UnJXpzTeQpwwt4/y7zYAVwxYzeO5cQuSDCdWQJl870sc/6TahNdKP10PiT
mrHq85RdNSPrCz5gc9YKqj4PfCb45bkTJd94fFy1JGoUBgQ680iC19dUXsVd1a5a3nLp5uIkVzN6
i1XBa4fk7V91Do0OX8fgB58oDSTD/D+YRzZ7CPp/AJfNFDoigs86wnSGFpDRgYeBg0+aFIFlLKGO
U/KdZ3gWsG7JOBCTtQHVtjhc7I4y2Bc05KNqh2ZQetSyvSFeTNUtHk5hKQNEZCT9rA+a2Q269Upt
kWF8hbGPo+jxjCXfXA4Q/NGWc9CPz1LHyVmaFCVuKWyDim2TVpLsE9GpgfP8s3ze+RLPpr2USKxn
1E9UoRwPBY5Qxha5+0OvInhNsKOYSsRwYGA4TYnpQipDkvBAYb62AaeVamm/j/vRXxqUQLILPW2H
nh1WrE+7WJt5GsniK2+3HECsqSez/o+7W/80sbNey5TOoknt/wHRGEKQzbqCIU/Vcu3nnfLgezV2
src9p7ev41pYsTRyS+qMfY8eDwkooxtFLop1xqJxD0mZwZZwiiG+9ZnzEQPEYWmKD9cbcSu2q2R1
PQsEXTKAJuMC5JsmvURScUYUsfKjWjd7addDfNnwb/fviWcH1RWB9ZQImw9J4utUNf14gJbstuyY
tkD6tZeUu4Oh6ecrAGG4bN1Lz7rhFI96JXbKgCSEIyKrXOxsfl4S5WQsl9WApXuoRjEpANo9SkFL
msS67pUxBZIwKllIsVTFMneMV7+EfHmJnQoM/wv0SwAfus1JbijKhSntLHWWPH4CfU4dbmj+5zuh
wYY5aUgpLSpHI7yHRz6cW7CiFLNDUll07/qukRdjXWdz6x9H+d8+878frikWmvH2vCvACID6Bx+f
qMgwiZWp7OVnxXe0Ro7OPPDixM0b7CS8y7WBdlff1jvOJSCIWXpZdHgLNN2gUkCTB54u+1efIIG8
FitBzw35ykrY4jI8kX4k19dXGM0cYhFjpewdPRda+OWn31YiS8vEE3lK2v/65E0AJlJ33SHPk+Nt
zSL3XZ0znzzGwi2hA69AaqeTWq9XE5TSmqkjpFQlOZqr6fr9H+lYI3ySpfR8iG4+6OPwHGuJ0Tvw
nBhhiX8w5ap69j78r2IDXcNTtmuTDHV1FCtHj9YV4hf1IFSQZ3h5oodhIMST9v68rLsOUKQBBd3E
72PfCJ0OuCNhqmghtFsB6tGw3kXg5hgt2aZApTxyucJmiuxRrMUBDEer1jkhQNNsNrUkwh/aZawo
tWFP6aBq95gWQQVB+vtXRg5AyxLa41Iypkvylyzkx+XuMk60nLMdQSMyjjFqSY7scS/P8CwoOnix
vEZ8X4V3ZOi/z5ooJic3iLAfZUOMrd0wh4Cm7GYCDQvOKUDTfFo9QHOHu4OX4xtUm9q9oOOJKqz4
JScAv4W6brm9z1GXQKnQx6FGAPtbJFTgyrk7ipD30BisrTpUwv0R9shpA6klZZr1FTXhv/ie7auD
kYf/9ZDbW1pLRl4e0Wt1QZuijpivu+WRwNQUIVZ6K4iJb4VVqY4hI+4+iQi1X+G50FAeh0RRoDjp
CxB48gcY4/uJUb4fplSjESJI0eq1PTHjQJ5zmoR/Ni9d3epvsGXsvpYImYCyrdOcNlzbU7I1FUWd
TwMBN6XBedjYDMMfJJX4dV63zV2IH1yS2ts3IW9lKzzpVwMMSNeeawFFCl2fVKOrSI1gCJK529A3
nPLjb7V/fuRZCoVzsMqNEdhtzRTbdEFk1YPk5RwfATTWZ6vojVqldVsJYGe0cuJnSAhVuq4CiGAX
XQlU2R4b7Y9xZrenaE828biIb82iZ5pO/4uLDhtFPg53y7yXwMJrJUJmnrODWxJrA+UNPuXAc/n2
PN737bOSsHCmLt5RRC1qTpBmthI8NNWivBX1kGbcuTU+5vIXa6BnfQ8zhJgmlicvWvMJBbXJ7gvG
MrigB9uuVJajHLCp/4545gvmus2KQ64ai3U9JznlTdZ9ix3m0qxtFj/euAr3heWtEpq+FXdgRcYl
Ie3jHjEOZ0K7FUC+8BbWwMlndSyd5dA3Av3P3TqlG6CfSaGLaX/PA4j+ENhrzmcg2CyozcPaBUs7
QSP2Bm7DnqVDcbf/5dYpvIXgwUq9g0WC4IqJLBh8ULFk1M/xrGgJig0xPYG/LvCk57oNTDH7E8JQ
SuadjP5mcrSp/FBo/AU54e/BLLkEVbi3k7wsHolWnAFcuDbQA0aVicRu5R2DJDpLM5nqYnHWeoqh
5I+l3aEvxCZzsVoWsQn2S/VhyM5Q/BMCgIuDeSz7I/pFq44ATPsrrXYxXMkFVYZzsjlEu6xzhTSA
DA4WVH+jlEUNGAFcaKbg2+Ge0Ulua2Wb3+GDAtFDUnqIekbDL8epjgTuBUK39mWnujrD6K3h6Ly0
l/vSTbEEUowfVslDXgkaMaPpFuBEXjbPg+0I2nofQ1V1Hd0hpkjvshkTn/OY8ZLbw4jb0dRV9yAq
XHvqYTtC5DmxgdK4k/GaYmYkv2h2cgDqXpMA7/i+jNlUwvuHKn7C8xbPy0lUBMSxNZjxWQOWx2oD
ARSiNprXDPhSywIvncIAljr0+UKYEyG8o+gYF5b1u6kx9tugkBGGpXuA0jsk4Q2JMvgM3eDLJFpo
ovx9KcnjGp/5SsDgpdmwrrfl2JfmOxHkj3/CaaQMk/Ukv5/93kGCvX+/daGBE97VThRBtG4D+sY1
lRl8rRsbDm7kmX5fevkNCmKPzCHVKry4aVr8+ZP4vLQTpuDbcbSZhs/ZP8UXum3BfYlk2pVm/rco
QKM+K4mgh0VnP8OUgcgMmpovulmcYJ2CZBfOCPHTeDaeaYMQfsWOJe2MI/Cg15V8BFdBDALuFYuo
m9l+xZoER5Y8mJkEw2y0SJVpIXNzToB9BffHZrU0XLMPVgVpqrbRCHBeqa9C8TM6o1uNulAV4dlX
IkcOTaL2zNzov9UIXcRgou9D2ocvZWlfFgCJ13CGJ692x9SrNnyWV3eFFOaZsxF3dKs85Vw5s1Mu
h9Cfh4/TW0RftwKQlKDTRrPSrt6/XNJN+e4A70qJ5LJZf0TmKycthLJXbZL51OMco6585J7LPV+D
yc7XDHSraArZW5hSVqOXMziu/Q5o3KHrYdfmMpKrY0kz4lnKBIvwAFGm9EWJBDwM0a7d5wnTcNe6
zYiYw7S+uaku25yMcI1ZDDLPXyfRJOCWJd7Xnx7Xxrp6APcVgI99LbDg094e86Z60UzV05QDWCcS
ucGTsQQ6VRP/Vw1/o+deQoJ/h1KUO0fB0IBRWUUrn/5qmf17+2FY+0tbbAyt1ss8KsiJSPDzEjM7
1+c3Km/kSS3fP1HMY+4AwJQcwwG4f/3AvGrSV4DlvYDunglqvSqGp3wahoqQ44Q/ysrHkoMr5d0+
mHKPOHODevciN5TkSEnO20iemjGq6L2shjOWHO7oQmJqyNz827Cd+MowHqTEyUmUnc/6GL1M4ZE4
2qnNCpC63cUuqjrtu9764bqbU6XHJuymitSZ/2EgrpW+8u/B72t2gM1eP/wezafBwThKaLT4IB3Q
VEr8mIOy6g7mAPZ/ee7jpkGOyA+RibFMjq8M3cy++rDpDM6HHv/Jfvq3Pq2VrMgpj6E5q2hUowO8
Ms2cfOh828LJoOsehxrEIUhhM5F2qbz5OzAyUrRUsCITQssUEIBHJPV67lcYoESaSxyLxe24jbRv
NzBPX3kQb0tahz2CGlQJffWJDmDwsyDEPKf3Ec8muxK527K+2hME9axDUMotYliSEbfZ5dUovrk7
Lm/N0Ylo2F8nT4Kf5p9qqlAhf2VWWC6bb4uBLD62jGNjKQNfC657t4VDn3/DAndTYGn260vBGHn7
bG7dS/JzetwT80BkFKKp756x+0QlMgHIzJ8FsYxhg8NGxrK/vs4NrLYiefDfXDTUVXyJUsLtWFPj
vgSum9TYFoYNk+k73dMoumqsAOhUNVqUw9oEpc6Ka9IIRMawHTacK+aZVzyR6JJzIKEKodaCLdAS
2Y4jh5uUf/HPFuZxLqZaCSyRtfoQO7mY+6HwrcEYVUc2C/Xg6epBDJaXvu72sFZEhRjMndpRXfoV
ohceJ/UOWER04J/5YVjZb4WGgRyYcbwlEMB8ARy5yAYLbbF58Eiwo55OlGDCvim1IqDQEtI4Wu0/
qDXRo18tblNHMBwFuYchExfytsbxV7qjx98zjIHWtSiUfIF/FD/unLhPQrFYoyUX6wVWc49URdBf
BJem9WB6alX1e5XxkrHLha1xKTEvnw5ACkJlKrL+nzgIARDIQoA4+zaYclZpa8Ir+pDCNorSnUJp
HMpqONY/KWxIacIgcpCcU0Ytsn8fvOcrS54bZSBHog0H5w0gt6dpEv1kKkgZx5fOkwgLJVV9pNb5
SqAl/Meyyszc2aWPo5PqMmFAEWiSEh8aAlfr/Aa5xLqrypeMpy7MvGqss4GNRqWKsQ50mlrpVoyY
VQkqCtes23DpN3ZmsNnQucYB1q4H+/v5ycxfQal5GnGgl4Dx7FrTH9APUPw1wsNzypKoA8ScX0BL
tFs6wDkuyeMkTgVbGb2LvQjYCwzF1HlFiuoO2QxD/kcs6z0DOlJaJ0HXD9jOetIBnzZLExA4kToj
umta1jDfkfrZkDou4ecZLGW89tGyeU3Yb0Ojg7X3Fn5qE+S95n703Z86wE+2jksK7dkS+T0gJEb8
nyiPvlZcszdowuHTo0lbQ6i7lsz5z6Rx1BbTqFGO3aYBOtqD5V94gK7Jm9RTG2iRJlPSEmTrHcnd
UuD0fEui4vw8n7sck6BrT5zNjUn6Eri+Vb7H7B7KPl+XpP2ubqUNnk1gXVaLxIkO3pUBPC31NqTT
BwXfevR1PLGefNXBRSJyfbF0aFMB3mhvSAlNdcrgKdvgfnM8nVv2gFf6jS/h1oW7/J8Q4vAvuWnG
rW04VtJyh/bQ4Ltew35s1i2t/vHpb5li66F0p17Mhz95GR3LDR9VPhCPZoGDkz8gbpcy1KsDOjpA
ot7gWD7DCbuLLhvy7kxj4QuTdnSpqUiIskaSPr1sibNPdMNeV7B8ctcodBlTCPN08iAj8B1FMk4u
9BkxzslV0V+Tx/n1vSwePDF1Hzioo0hQAt4CdzhatJzekWaPKUg/j//jJcU447ibRTOpViMoLiHo
9FrMSfZ0UgwNGYHwieMTX0v+6i7NO80alDpxg9znS+2cLMopJqWKIwplYkI2F+dI8c5l7w/hby+N
2PxdotFWgOpR5c+ieBwNLpxd2Sdida1Fs1h7eUL3f38Au1zmXonfxUyLG0r0/o7N3zrdmQlakzVB
ROwmJc2+MIk7wEr5ARSA6iDb+QD4bbjDIeniSLyMyoDmVnmkiGD80lF6r5BYOYetKTLFj+vJVVdr
3ucj1bjHov8wdJIrOGJwlt/e65SwAgiwhRaroTNvpCa6/xoOb0xUqSv94R0sCc8SPw1eaXE1ZrFC
15Uqym67UT3QMO11dMG/lwtDL+icQZ1NOvQX31VeNrQlzjjC7AlNinAHDJy6bEHxwPNVFelCCgab
gUlWUQ65M7waVx0hFiZ+oiGpt5SSlHb6Qgegh77rneNVH2K6RMxoaHKd+NG9Uj47SQZxeVz6Qx/c
kK+ntk990C6FTcgr9QlwoyztE70YsKCi4x2PWTAbYngMGWipOJX3AiFAqyl5hyUJUjbWB0BYuLUV
WyQppzDGkm0xKzwG87zjNcZS47ZygtStzYqnoBc/ouJVBDO4gC3i7LCX+h4iOmtJ471gFvDVW/0n
098ws9sM/NU6Up+MVNHBxeUSrpTKl10hUbs8VLQCuJg2ythBNts0KWpu2ZUeQ30vMkhKkxJhpYkJ
hkHfFxMVr8LA6EsI+nc7xqYykR64wgP4tdirpNczgx2y/Dtoh8juDNbxpHK3EQ72eqxZ1+NR/532
/QQRxO1tVCLaK/SK29pmLhVOYJZ9m+CvxbatFFaezbp748SWcuBUPXdOLBX5ZJevAQWN6Ex+WmCz
yQnSaGhFDfoBPZLWky4WlA89lJWvHoE2rpAIKR+RsFC2VbLo/5sagT/vLdKAxH4cJSf7AOp9Km1A
WFb9G4pQHDKS+GjwzH+37DcihFjVsJ/3wdYIWo7U/R843cAirb+9qRyYysNlRN0fmQvkUH5NNARJ
nHitdb+fJe/IdDRzaFVz3z4n5LR3WKtxVMWR25lgXWXTUWkcKpTwRgGIQ4VaUYh73QiqJFa/MMWh
/yZDkwq+gr3Dth7JWkwEqTJ3LysIb5lWTmivk1GKCy3iuHm1e8M/hbGA0B73HRdnG4CvKO65xKzd
BkBTbFM+Q2x7ezzjyFORHt/lMmftt8HkpGHj9lHr0yyAEcIZt/E7mmD54a5gcDlaK0oM3h4vkOkv
pxHt1skkMAdn5D1JS9FXeclhHHemKGrH2idPt5N+sVjmViIqq50krlMieZ7b7Th7AJ7d/MNb61Rm
edkQ+dB1NenTBfi8j8kUA+GGG58kDvXgNGNHBycOJJxXomqHsmnCqofIIrWH45t/YqyFC317PsOD
AtpTns7Gme9jDZfx1tbuhVC0nS0gCS4KVm4sWYbku3i+N8C/X3mghrOdh12LHRi9PkIKTaNWt4Bc
emxz2IwcDG2su9M+PG4YQ4BDDFS88sNUhH0oBY6UphNeSqqifoACg82gQ+plScHo46vw0/W82FDU
hMlGcnz45r9EYSPz6zjlyieRJUvY8r6ai9GA7lswnoU+j6c/WaAKdKioIuQx9/IAKaDzLaExs90k
f/NOMNMIHqfhowOgCIRPjxGj0mmftEopoGk3wXlRI3rZ8Gqt8RlFuhX4y++u5ZToSoITSDpI8xOl
rml5WnR4XpVO6cvnEaLnkjT3hJnoXnsmXCTU6mDmveB6Vph7LodNhhr3wlKFLg6J7IIR67UCtILs
olNQUn+cr3DTHkT+kTlexgYYKWkDbkC6dk7adJ/Tq+9vvaONKExTERRUkThT6ilEAIzdztkjmRn9
0D7coYOFVB2o/fWFocDa5kwRtQhK7Zsw
`pragma protect end_protected
