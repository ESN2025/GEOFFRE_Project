��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:�1A��"iOWV��Q����u=}-w8��-�� �̠M�s��:�Q�� ���Y�����A���w��PN���*���.T�����Po;X
1���8��Dq��?�Q-�'���g��:��Z ��� ��5���DY�9�ҿ�bӦ$�l@+�mXe����1���-Ud���ӷ�@]"�A��|&WC/��6Wt�̩��V�u�H8pd�ћ���p�/^/��3�}���jsc��]!l�%��E�+�|���DD�zk�5���Qr-(�1�g�+P$o��nTM���E�hN�j
��N�'���G��4���n�*�aK������� ��s�	���A"����	m��8�f��dJ�K՞�2���Z�Y��N���T4ŉ�LV�2wx/�:m�&�=�9G�=\�P�:)��߲����C�pR����C�͎���4O!G���J�BL_M��+���o�yY�J����-j��nBO8���x�������<ģ�ϭ��+X��NWo���T9��O�����
���'3��*p�yE�^���e���C�|����Z�%���	L��9u��fC�mWY�7W��[J;U��J>$�g����|�[z�3���ȱ�����)��^N�p&�ݦ�c!E�mj�HL'���X�zl�	��Ĥ�,�A\��4��G��C����r�V�vi�NH����(������⋵[�(�R��v������`x�v� S���㞈1	}�L�N�g,���N@�vM�׬��R��o�T��[;-�_;~z�n�P�!=ݾIG�R��ﻴ&s�V�C,�@ht'��<�(&Mn�>�'�����Zy0R\M�n[F|_�q�_
7G�3�������cf[ݢ|��%�����Ռ\[�wV胟��LG6���3�n��J���5��	��{��h��AlU�6��[�ʑ''*ǐ��&����e�I����|c��z�nɈ��C�S��)|߼9���홑v��3�c1Cmt�'�(�ɧk���r�lR+�0��v�hq$`Eq3� {�=�+{a�M<�kjʮ�Ѡ+8y��~��3O��6��RƎ��.�"���ʖ�>�fͫ��$m���KL��\��޺�u��|?Y:�k�af-09 ���̓��HÒ`Û#C�"��gig~>J1��I_ٶ��,�=GYwO%�ˆt4�%�� ��RkR��}^�zϤI�� 0��q�3z66Y�b޷.b��2��V���c,��-��M�-�9,�F�F}�`��:xQ���*�ܺ'��	��Q�HN�m�z��h؋�ip��75Z�]E��������}̢�羋���)�gV�@.h	�_����=��RO��ՌcZ`�X��
e	,��[���#���f�\:9R�"+s��L
 h�K���P����i�� ��9�$�]ctRw��cRn؞�T�8��Q��ٔ��܎�J+䀾���:yo��^L�P05��5a��(�%U�X(���K6Bi��'����4��"����@��C��^6��u�7�n��F�?��F������y�z<���c��9h H�<���r���A��.f�H����4�I!�v��X�&5xeSX�n�1y�7,% ���b�Yf���ʓ0��E7��,�R=����N�8ڤ��)�8d�b��wSdWL��X�H�p*m���Z�}���JY�/����.��-�=�g>9�OCO;�asӇx���R�GET���YT���.�$Z�Q����!4F��ߎH���F6�C+��ׅ#��3J5q%�>���.۷R��ڜmKR�R�a�CQa(M��R�TD���NJ\CF�m	��[�����2Z�cᗗ��'�?��FN�`��\޼�s1!W�^����Bew�C�z�I����w^���c��NK���enc�˻��)e�����E�xqi���T�vtV��QB�dz�?�t&��~<��y�s �"͕Rk�1�{C"��P� ���ǈ�3i,�{%S9p���3�h�6Ʒ�VW!~C#V�n� �NZe��)AE���Bc��X�0��l�Zd�y[7�x�h��ܕ�QU�M�/���Zg��7l$�N?��hY_�x��b�FV��#�(�,�� �3?ܭ�ث
�h��;{xE��)���]�Ѡ��$���0���������s�8g���K��<Ne"�M������ ~����c�(0h
���[��%���;��~�N��X��CM�{�q[��Цb`R�s���� E�B�f��M����Tc<�lv�0Kr�v�����ǥ �/�Os:ٞ��ul�-"�<�
�x]s�&��i��͸�Ʉ^ a���s'�C����ɓ���V
]9}|(�+N<ь:�jF�T6�	�Av���s��~����n\[��\����������Pc�Ѧ�~�����)�����^�u�7>���|y}<1;	Ӟ�Xv@ɗ�,��)�������6� R�a7�{.��O&�H�ݜ�wQ�]S
�u��^���#�>�R2=<�8wb�I<�,}����]�h��:Kt����-��u{S��v؏.e,w���/1x�M��C$ueƨ -� sւ�IA�[��N-
��_��^�<�F4�Z�/t_��-x�CR�k���QR�q[k�@B�uV�x_#����|Í5($���`)��M���Np`ʚ>	F�=�Ysf���kh����K_�V�t(�>�7}��&�j�Ǽ���h8s��̃��m��'r��+6+1 ���m�[�����w�3�Hf�,_R�s	#`b�9W�/��]���M��c�W��B�$��t��Ҋ(�c�o��I��/�`YK�&U���$\��J�aAQ�]��;B�c�ڒ��|��2.�.�1�BZ�����3���K�?�M݁49�
zu�	T�I��J���d%�ň���p�-����B\Cɱl���F��`�]�`w�;G7X���R�ύ���eyP�j�Y>�0�ݿ��6��̰n%�&`0����s�D���	x��ilD��i�o=�:���s ?с1�zNa�cL�����b���	���f�~�(#YP�q?|w���\��r�g�,��)�����=�J��G�:�#vs�;@��_���O�6��|>c!.�1�8zJ��~W�RsR�ͨ���V}���� J� #���=���VI�=s&��Ԥ�p�ÖkEp�9�-&�>BΦ6)��]1QJ�흳�B�ԒPQF���t�Y�|�!6�w��#=�2�38I9�[��,�����N�bc�Dʺ����o�*=���om�O�r��&���4>��@Q�x)���Q�B�&�
M�Zv�L���O�t��[
�ɞ��\<���ȑ��D�'+ ]�;���39:
��A:�� �kv�ʞ�K���_���2�u6���q�[) 58�S��2����O&�h�����|��wν���$���0��Rn��lN��0��ǘ�Չo���ti�hΛ�iS4�.�8վ�a�M0&s"۫�����j��
}�m���]$3�b��������J6�=��b��?L������қ�x�{x?�-H��_�J�9G�w^�%Đb��bn6�Œ������%ʗ2�~�I0��i����j����Yn�7h{C`8Z�I.mNb���,��`4��
���o7ҧv<��`�'����K��XrR i�!��N~����Z������Z�6� MJ��/�$OQ�|����-�ee�KD�Ş��_�ϣ��������n��.�~J��Ii�􅜧¹k?U7X����%�uH��ݹFzZA����U{������	H�	5�]7Dw9�x˝U���k4�S&X�(k���2���`=]\5iL���zx���搟x�<��pљK��'�fz�z��9<��ϻ!�O�^�L/��lh�x�z�%�~�ڏCz�L��7D%$���q��cE��w �A��4�Y���El���b��肓FP�>;3�	K���e"�s�������%>�ĝ;k���`r�64�j��S�e�ME���Q�<���A��ańz�����Z�hn3w��'���]>2잓�ۧt~��@�[c�ؖ��h
��`�2b�p������*Ň�E��>,H�=ZwҀ�'���{�*�b�[7��ĝX�le�a|������9e��$Gzw�����ٮ��r�P���a鱳7��ZDm��@�\���r�o�v�6�(hhA0�r��ݦ*��EI��fo�3��|1`�x8UPB���ޠ�0��Xv�Zqg��Vm}�#��<�1 �f$�+����ۮ.@�1�n�j��w`u72�~�-���h�k�Ӂ�H��~u�bd� �V��^��ѿU�R-+5^���>@�ms:�!
a��G%�w�\!�QZ0Q����;Ԁ�����=��uW3��f)� ��^�{�U���y�Z�����^,�y��>��m�FE��������$½fo�*s{[�ѓ&��[A]S��|\����ق5.�fN�J_
��L��Ţ�D�nș�:L" >��N�%
�jI|��v)�	9@M�+<��>��6��'qQ$���c�#���-4r��"�hHS��0L<��ٺ�*�F�V3to�����(u����X��T���~_P�b����c�l�~T�1���
`�Y<"Y����i�lH\'j�Ɠ��0[�X������i���52	��:�0�Щ���։{
��z3��%B �5])�s��0wa_J/\8<je�'ޘ�.��Ǳ+(̿I�Nb>�m���(�;5�-6~���j���G��$,�����LP�c*T��p�%�y���r��y��K2A��������Gˆ��f\D>I+9���p���n׼uÃ��������Ȕ��
i�m��lN������ܓ>5��Wt��(�����6�����#�b���O��h��h%��G�qH �y�v\�!4d��I���m�9���j����*�'�F�����2q�O�	Te����~�P�uR6L�99��NRG�N� �]�lz%��aT��Mu����T�/��#\Pb���>�,sFf�(�`'��}���y��8�6���G|䶁��Δ*��
�5$��J�Ɛx�Z��c}5K��k�N����^�>VST V7J�[�.4�C�/�ӳ��K��w��¿��Y��%Q�0/�� ���AI��͉<��E���
����w{x��\�@�bof�i*QK���]	#������ET��Z���#�ϭ�K�sF����}r�l#��l��94����'ٹ�����(ߍ�^X��k�ͮs��v�3tɿ���zx��^�cj4��g�Z�V	�&�3�s4������S.nl0p���
+���v>��8�V�Ut{���$�3�ew�
d�k��6�>yQA�K]�{�<nh%�[���	0�=�ߋ
�{=��iX�><@���1�� AXux�6�3i�'�s�K�a�
/.H
k�����+���,ȕ/E[㾃��>��I��ä���3���3.�7h�k�{ETmoJ�s:k�z?�Su)��u,X>��x����\��һ��$�W�2���+}��������Xv�לm��R������+�cA�^�����c����ߴ������*M��<�HU�qq���}K����3��;�(�K⴩�O�p�ހ��5T�d�Cƻ���]Vl+x)��x����E�2#�	h�������\aٱ�/�OCuʝrŽ)�z޴]n��m�2�?wMެO�J{�:��u��L��_�䇚�i�ђ��50#Ie(�ϒ�(�����l�͘���lE�>�u�/Ƚ���	+���B�;�z=�"��1�II����
«�})H�Q�R�c�h�XW�㽼~@ �߬���nuS6j�.�z��r[�"
��;�q��(L���_}��|�Z�Q�X�o��Zyt��2��$� ���̛ ���p��/���'�{?����>�'K��4}��ȄW_��7�q��P���Ӝ3(��N@��,�W�O� �
���M��Ps�=�G���9�`eo��j�|)f��%|`+56�.����X.a\Y5,	|>~�#����T	���O`�N�i���R3��D���LQ���[vC���R�O��8��;Vq9P}N�b�wB�����n��헞��̣���#.���f��|1RЭ���}\���_��D���3�� �Xo���1P��PF7�-d����	ݶ��bL8ڂ/΂�E3^<�5�E�J�EЙ�z���<^���td�U8%gc�F.�1\ZG�zE��ߌ<h|�z|�vB�6t��G�yN��a�'���(�i��T�,�}Q�/Ө��3����opT�:�c��.���(�uУV![�d��Zʚ%Iɋ��e��D�ӻ|��B3����A8�ҚzA��H)�{/g�L��9"��X5m?�BΨ�b�Қ�JDjC�/b�?���������>�{C��٥d,�����V��B5_@4��T�6�b*ӻ����B�Z{�B��Bv3%��y\o�Dd4���d��K_��Ht��PJ�S]*=som�]w��Y�2�1�w���VR>�~"��Ȉ�N�$[v����7����1<��4��,��:�o�S�
����GjGE�2%L�px.o_�
x끡����eݓ�H��Fk��s�f���b,���J�v$��Q����X�ʌ��юy��_ڣ�J�4%"v+ٽ)ՏyJ��@_W�U�S���k�"�@��u�m<��ɗE8�A���|�W��pG�7< ���?U�dP]�۽���\6�\���$Mr�T���4��缫�)�I�`%�2I��v�qȌ��B�����p�k���Q�F4�M�BNnTʛ� �}m.��2X�B��y�TI��E��?�`�"��J_���iՕ���P���9��4|��L&�|��w��q-�X�f��A}���h�4D ���,	�4���ȯq4���cq��,	F$�;H5R?4�}���W(��^��'�^�X���R�_��n��]�z(�r�J�-+;�&���M��E�5D�\�L%f� +��s��`�.�$V��r�V�Z�Ao)���G��Vˬ��&�  ^����PW��5Y������x�}��sC`9ٕʾH#�i�T!CSM-:E���]U���-3�%X,k��6/��ʿ���aE��]�/��0��B���J��籩�u�yh8g���@�����������ԘQ9���+���.8gW{�Dm�ؠ(�$>īSA�H���.�b�wK��4,�^v{yNr<ӥ�4)ql�[s��#��Կ��4�	ɼ�tQ1#̶�QI��MޗyIH��<�Vt�(�?\�-sZ��1��FĶ��n�!�-5�1�c}��O��w����U���0�J���R���Qк%�o%˷�CR'��	���x/z���%�`F�A�];ON��*��k)� �h�.1���?���P�)�3��� �vX�c��[�x��r�.�׌p�%�A�!#@WWX�Z�x��G�)�z����Ȳ��,F���Cݙ;���F��~���ď�T>��1c�)=1A���đqAT��|�@-�L�j��^ �V�7��!��aͦ���z� �#٭֣����@�"gDL�W��P΃��#ƽ'�E:�����/=��f��z�[�+���ʽ_�x�^�"��>J-xwWm�=�&�O�G��|ˍfUu��nᡴG��=�8t�42����O���,zN��~��T�tR�zN>�7aN@�R�iM/9��r�ÿg�;ζ�a���$���q��jS��T����\�H��L��f����i�*ne���Uʹ��`�j�щ57��� I$����C U<�b[z�����S���('k��#R�@��t1K����6��L��z�Z�/~���V�"}�i��PN�Г�޳�ہ���A��&��C�	΅�f�����uN�ܞ�ڮ��}M̃b�[�p')!_;�fo�)��#��s�H��1��J�"�j���Q��
J�S���8��M��� >T��9+ӗ�
\S�N)E3���R��'�2sn�˦��;���)e",�f�&�'�{��"2� Zd���Y^��f˕J!O��`�� �!��>��Q3j��P���3��e\ �� �t�Z��*�"�^�<���p���C@�m��r-�l�O#�I�k���B�;��&OyQ��q�RR|^z��@d  C�ц*क��b��l��������ţM	�n�)=�W�c��Ĭ\��y䌢�b���S��a�l���i���?�5�A�8�q���.����a\���lvC��S+�&#�����i͙�c���O��M�9)���#�83L+�_(x�"8�Y����T���Z?-�	�.;�i6?W�"W�(a*�\{�:�|�hda53;��vb��}� �+���@A�\���L��>P�sY*��{�(|�Z%?(>(�؄r�V��+�'c�ԓyq3o��N�$b�XM����+��'?x�;��雓��+�WW�OWCD`�����V�({z�T8����jG%�Q�g�dy����t��^_;g^��>�h��>Õ~��O���[�_@C�e0$�8.�/5wHF���~ԇg��Ć4�|�N޿He��Č�Dt�
����蜓��Yx��$I�����%me��(�����I�ɯ0�̋����[ɷ��:e�K�LυE�u��4��E7�DEL�%7.���ffׯ���7�D�I�b:i��  v�H��y�C�T�� tf���e�K��&�5��uC�!�9o�&�6Ox�`8H�9Ҹlh�m�<����\m`��v&���B#�����y��[�2���,��K�N��,�\�3؞��mE��"�Z�:�Ej�O����\Q�F?9v�O7�
M'9�/�ݾ>xi��GLd4�|�bR�ua�N�q�����R�*�{Jph�[u麗j�r�F�
Q�Ɔ�@�3���5<�Z_G�Qw�p�(>x�	G�Y�_�U\- ���2Ѯ��M�!�Y�U��Ye�5	�l�j@?��v�(C��Թ�͌{WwT�-��8�.aQ�ĵA�-�O@��E4����ؔ�ڟt�顛��Hh�����/?<�v�!?��o"/Hl����Só�f�$���HT�X�%ͼ�l��$��c�q����V��p��FO��Y~�.L�����8�g&�j/���xA�J����>yvH�L`�J-9F�@D��d/8�I��Ě����r3����_���{���*�2��):��^�L��kJ��=�X]��T��rN ����s�%�� s3�b�vI4b�[�r<��H�H�^�9�2 �Dh�wC�v��M��|�H�.���{���0�.5ט]�K:�!�;�ST�_9M��U���
F�E(Y&��9�QLЌ����B�>T@ū��	Q���/y�8����!�	�gy��8���p���x���8"I[HR�lq>w����3�{Ϫ���O��*j���56$[<-vE�7f�z�b4��,�-�����Iťb�P�ٕ��B|�Պԭs��:}k{
5v_���T�
����:{>�8�e
����|i42D,g��1�_����x-�Nr�32|
��������e&ͩ����+R����}I�6����߽a~�l+v5j:�a Q�h����a�N�^�U%�6(��BZ�âB&e���n�-ѓd�����).I[J�W)e���6��F������ñ�3��\`4 ʪ�P�uV��������Ў���5<�lXߘɂ_pҔ�C[�4}�
�q��!��w���GsI"��ɡ�[o��N%S���!cj�~̷�q�o�Y�3��d����ig�?_ _nQn��JJ�I�8J�z�bB=G����dj���5���e��X�
>��S�ܸ����Zfr^�ꑅC�(��A����`��\����$�N>��o�j�yϡ�^d���<�<"ҽ�|:���2�P���H��祎\�22>����k��@(J���T �-���&���ܩ5��,�&6e�]V��1]�e��_5"h
@�G�#�r��ƿ���*Or˦2O�'���.;�#��p�����egL��������ş��xG�S������
|{�Y��A{k�R������icU~��.�i!:�m�(@�i�
$�b�d6TM�;��2a��\�g(�,�����%�Lо*�I��R��4|���t�'�S�P� V�J[�>f�����_I�}!�I}1��g�ڙ>3E׫2�2kq����ͽ�sy�a��A@��.���s&�q�, �HH�9���0�E,�Ɓ�Sk����x����f���[ ��Q|�+���ޢz�?�T�g �H�g�K��P��}{�m��,I%����)�.C�2�{)��$Iڶb��I$S/�e��1����Oz�����@!���(q�q�"rr�:�:~�����x�T��)ZT@���ثh�ZuB����d�7d����}�����fx�j��M����t$3�(�)�{��)�͐T�ڻ�@!rz'`���� �Q���&�?�g�Ҫ����-K�)��ů�f����M�9o��M����]1'M$G����c;�q�z� �.ڵx�v�]s�	���IT�}ň9�=ģ	�_)&@5K�Uj�ؿ�0i�%�
]��˨˚�l��q�tg��+S�g�Q6�a5��k�>� g�����Gɼf�~� G7� ��Q�2vL��U�a�d���g�ݲEV�������'��EZu�v���	߄�M�4+
kօ⦗��w&�P��]Z���+&ă�ZB!*�c�&��u?�@�����E�+/Q53����>��H�}��/��s�8�5"��Z���M��!��L��l�NS;wD�
�3���8I*��ȴ8�	��Dp����
&��}ȭf6��);]��y��N7�'@����W&��>"|��GU����;��,���%r�K�F`f�>���)��k���ۀ�qL����jZX7��F힠�-1(�2(
��]�J�U���囖}9y�C�c)�v61����F�>�������sޟ\�P�0���`El�=�	^mZ:�c*n�l�O����	�>�!+�M/G]���q]_��4��.�+��[��U�k�i�+��.�"��2ub8~>��`��j��S����#�=���8Ң��߯�t7s7�r���{o^��AV�����-���`���JQ\:�\M��ؓ�n���U��}F���2��E�6ڥo����[ܩ���>�JM��>n�!߲n��T؊����H���o�?��'O$��w߱:ME��q�t�<�#bR%���f7��faH��/�|�%����ٟKu�4��j���� ܜ<�=L�d�Jp��mԇ[7^����Z�4�ы�]������L�I"��f�T$%[�1�b�����w���z�K��I]͚��E�^ܪ��R��Ahԏ�rfTş���ܴ�_R9y����4��?