// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:26:03 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MltU7i1FhwTpFzdSUE2voxXs35u4tnOUYqyUhc32Pz476wZdxNjmTtbWlmdVDARB
5uYYIHujwjoDaEbn/f0phdukxdeIVyBISI76OoAvR7tLQYqZgTMsPQS8oPHOOCX9
+REGo2EaohwGZC0XIp53JOpmckbjKmmq/X2hZfGYkd8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31632)
0yi6irxMdK8zmOs465uCCIZ8c87s0TOX1w5/tmsL1QWX80PeaDdhCuKlJr8lum32
dhqp+MBT7R4SAnVQLiQjYkArvWoZLFMDwewW4L+AHyz4ZYcaR2maEcNnT4xiOJ7+
kp3xBLxRxkFV/VqwGOAJHODu0ISZnMDucil3B3VawM3bbWHEXzjcywcqyZK5n+o1
+q1BCjwI8b3A+aG0+Z7lPbhzHZ4ZEGBGfm6HOyL3K0JmaojA2grHAqci8gF9zBPV
+sATAvpnJgGpbFw8NofIF/qEB9UjUH2RqZsJLy+RG8hh9l/Jl6LuUzjO94srZvbq
Q70vw6cnKNXsLKnfQJMN19wB8P9ODXPvpZAkAodtXAaIwf6s+xKWflYmOW2Q/oAH
/XtFOjF+pkFpiUFpcFRqXoNUOvUvL+uZv6VpYK9dWQ9huTX7NO01KDkLtvh5FLzd
Q0t3bbiQywVpQn5jfeiJwelW0cHM/xEAAhCAqrxJJZ+J2kdIzLVKlscq1WHKu8xG
h7pznjAnOzZpQGLyafv+x2gAKZNoqwQD5uBi3IayRFWl1jZGd6avQp7HoMn3cx1B
v6zTMn43VXx00RFEA3Fbwj75LIzfFf4NsjOZXeWVgQpLXsRZqYGjXc7ymb6SXZ7e
7P/hibWbNS4J1tSf9AMKZ6EYBK5KX2Dd+pREPQc6YsKJrPcdK9XmQtr7AWTFgORF
DR8wXXcfX++MAVaL/bQy7Riizlveeqglq3mC/bgUCdwOwraYakRS+UQN1TGBYZMX
sfAshSPC2+b3Vqrcn6xhrumhWPExdr6+2LAPn0u/dTXHTVSslfMEOpBArwrpbADU
YNLhahMj8j6bIw6ivO0dUhDmKYfM1GY2bPccjADi3krTBYIamJxI85Vu91knhbbk
4eMyM920hvCP37pPwX69zLlmyPegTwdobsV4cd0C/fuxT2wqMXlpSvi+HknoYZCW
eDD7Aceb5u4gGBUvrKGSXn2NMC+Vbyy2udk9fNSbHvEO/exhAXGRwtDX6U3a9LR+
U/rI+o5dHiOV/jszDVEOtkX/VHnXIVEAmki3JJ9UMskyOAWSRNaR9azmnZ73kfjM
FWCoYzXoPuW+r/UIy1PS7JhjYNpaEnqZmH+6hqrN8NobEdyz/5hweequ1SlHQiV3
MP4x33NPjdYfhBJokErpXiOKdQ1o3V0uQSc2g91EG645zwUzNW9aaCTUwS555QYu
rWIhyInDRqoaBR3LeGv+EnKBKYvzVMagfhKMq1KExuDWYFGYrRzv0ortZzWoz+vo
vJwsCEgBhX7skho2HoAiHdsb9JyKYwdn53bGe6pxSAsmc0lWuN2igupX+CaEaHvn
+TblGB8PPI3B5/Exr3W6PYURbd5U7Pc/BB0dwgxhG8cxPg4nDc4z0rzPYrMEpdIS
tkFQz6MKkqFb3yICKZ+uQNfpB+ANIKrXX9gOZv95RTz6gK6KSkv3MTAY5bivi/VR
EMLOA+MgMYODjSl/ZykKhRU2i5JW3y1Vc+i2ENl9B1dXRW/+gtRcLrffzFbT1HOs
cN27gcT8z5JwldyPWdsGi0fgvWG9moZz3G0AyR72Rpto3Q1COhWdqOaTd5UFT8in
XlYgzuZMbubDhDIFPpU6MalX7/AN9f1/nFT4O8cIW7X3iMsPocoZFnyE30KFgzuT
j+KJ+FlzZKBz4nFIJjJbHalGO4cLH9tG4Ug07S+ms5kNFEvIr/jmQtblVsC34FZf
c04FPLp8udsGXEP9q5VwCbxlrfzmHinIJopcKXtIMmXYCP9ecUxqBfeH9yxYeuwn
9eDd1eza5SJwuIlKo2wh/yd6/36L2KQvDw/s8XkWV7LPB5oGwe+wt/58NYPzjSfH
gufKc/7/ALFhcTzGzB7D/0RENjONATwbSnHSG7mwO7ed0xxVKywsvh8qP2imd1tk
WTKXuh9CWDCV4fufflxrKBUwT4dnvv/t4BtYrqM6e1Qud5qvPUWW5BYVYljdSuYO
+Sg3X3CYCOylfpujHhwrgk6cUUQGDanijkaOVr5EhAkC6Gq0CPtazqIk229iy8Qp
Fot+5+gpMoZmljDGxeSsLI8pzLSeXn+oPmHuLVsH9L9FtxWwWj1asAO+UTUHfQhA
K7wNl86qOeYqbFDvkC/nJPuppqL8vdmswZZyKvtF3udeRlwQbnV1RUbH1x5VTNR+
YEJj7qdkELHUFdOObizgqQ9e33lkOf921FivUOE46v8IMILo9yCV+Uzxz8dMAtDJ
1Zg3PwfO2eA020fn2Zu5UJHLLXZnexStqZj8wyRC9z3OgQhYPGihDf/QMGGNbljA
3aIRQThBWbe4QfrcToDAQhQrnfkI8rWqr1QbKFAK7n0Zn8BoHXnAxVtrL6dSTQ39
TaUVx6T09cn1PcUCvF81lWO1RZs7xc0tuLbUUDGrBXRjwBmL59gKRgtq9pQZixCD
XOO8snVHrXZJy5/iecsz4kuDxXT3Q97tbWi06cGCUiKxQ4Ow182dPdQGaSepP9Kt
Xfu12a7tIwHUCosPUHl85QVjmfduT4ACKEQTzEXfXy9OuXDpxRRL8of1LTkV/9+5
qURU8Vj7M7A3rBLUALGPDuBjQx5uM7dfKHlhK9AbK/nIMD7R+yWRwDAjo+cM/Oyc
/b8eIdV12IN6SNbPRhSaEtryHtQNn3zTpPSXh3byiHuemBgNs0LjPVXqw4NUWCvQ
mt7FqyFvjXJ8WjTKIw3uOKzAy7Eb0TJnrIifAwuzbEDOhLfwvokAwFRdPXuYS6q7
rgOCRxDVepOsPBRE2d0J2wiKE3thmedPqmTSsH5nBrtkj3qphZESdOinGTpFuPUp
djbvKgxhMGFns7pGT6f+9Nub59HUD+TMN4ssSN59Sk5wy33JoTtv3cI8loYy7nMk
Er2ONsjRYr5Lm3NVR+vJbxu3jT0nB0ChHa0+Mgb+Cyz9SzA2Su6cBoWQu1mRqN5Q
IBSS8Q6h6iynKBqdaRWTdp5gmL9d9qN2StSpPOefUf1jeCTdhPsDc00ZfCGkd1i9
dW+SxUIqXAPDbCDpBSfNHouLc8C+xiSS+mbmSELSEOmwn5Xfm8u4K5o4ROOY0x4/
vgCBU+wpFoxCVpVPL99SmZjtq/6FKLeN+ialnxSuvuRNF3AYrJ6d3FrMCp2x0tHX
slux+PcP4bC6bx6QImmri7gTO/HZ9IByGM41OyJnIHy8nQYsCSKPXYfiLM/RFi2V
47kGDiTQhakh7fAqJAasMmsbKlfKUGbtIJ4cw6Tqj78u5QHixLgaLPLIagGryQ4y
2jeN7Vy5Og+HvRLPBO669urcTkh9YpwFjDyFPHSlUktQghX1wXn4DyFjxLbUceaD
FAczr63PO8eovEvq7sF3+oghpiGMiLg6UnSSumBO/atagq0A+E7zXtI8ApPxc7wa
zpyonEZqOwbKxAriEXcxErwPMoh7qCqrvnyI8NENJzNCt0+5C5HKgGvOb1ZCoE1+
VdB/A3LJNLnT7yKBZIN1k2eN3oXZp1iFH8hf8PQjxNnZkX0LCho9b/a/XPmbsGX7
YqejvloY1prPO3zlTh1UJmQfIpzrOp47DDqEwCKHlc9riw8DUS+7kZJv0MRgmPnw
Tw3ZSsyiDRudII0lXwpzbFeW2R2ZIGZLDeRQF/HO/zl2eoL0kEC1kwbeCM1rrjAj
EzBZZ4p+nSq/sTWWc001lDU25pN15wQCJzqw/4DnOxGx4LLc8rNlrfVpk7a4+W1w
xmkIuit6sqCTS3KCyz1marDgTGPuVrK0CP0xIgp7z5Bz5Qj0jA1klM1dav5Sv0hW
2DhqrKM5AfXGFmQpepPAsnKvNckLSduYGckIen9YuH2SVdDVWUqXgO8repJ0mJwN
tXTO1Zv1vGfqE/Qf6go9LTSpa6XC6RGUVmJGwz6S7bNURgJeEIcl+z43TsnFp4vg
ic1oh6JfHHrTeii5kTflxR2CUul+XwiyeW0JQ7x1E2Rzpe8WWLyCX9X9YbBN32W0
hmn8DgEAHmyWatOFUAecJX8XCkFrZXYSFOXQLY8kTKk5qiQDS/r6xwciYFnwsX7e
UKbDlxg6fP1psOcrRxuctfrDkl3sAJ1m7yAyDHOncpPbS1cJ1BZgLEE+NiN8cKsD
vldV4v2Os59R8+MB2s/mUBjVxz0D6uPDS7SnpwL9B75KkwfBVvUdr/GK7RA3qE43
LgXnPkl+nxHTvw2EpjB8l3haILYCBUBa4HBhWdWbBpmcctITact0tT1+il3KHtK/
zXXve91KXV22xNvfIyMXzf+gVOoWXeXrEL13ROTcXKLv5InmoTiHS622EWBxYr7S
vtJkxRLUnwKNW/b6UzhUguKRtgnNy8qyWtxoP2Gk7yJ4WhFlTYadtAd7YDWLOFxw
dC46r93jN7afnHS/htnJxOKayP8AOp0+FWiKfnR+DfRIxD4tlP/ikhxrNYwV5mnF
8br1PPn7frqbmb8C+2xz/CzfHy/cIzr8uQnrKYQ3/IjjuwkBB2k/q/JnSjQmm/Bp
DX3LWK4d5uPqNX1XXknUB1vs5gqDljb8+G+D/3hPBWjrIhLSIoajtCH+qmFNyJBd
yqNIYRbYimjCf+CyI3fe5nbZLCEdh4OZ9c06ynMn8akbxzqA/cfC86aA+ypUqdNn
eo44vRkKFBEE5f0xpIXg5foo5crd37eWGCTY17x+w8Qd8yq3fKtXTd0M2nMATDZS
Nn0/+4+QTX922WrnQpg3z/uohYHSdb0MMTZAU563kK9muHLsDwtkLG7mmmqcckc4
KN3vFcMdkzMGYzeZyHOTWaHxPowCp/GTQF+An5mjUc12AbHJeCY2u3IcLq9lX0sK
a2dyA3WzAjLTZ0dUYPs+ajMpHJQk5KwJXymzcNJWt66rHCwWzwuJxedvZTJTtfdk
v0pqO/AcJaVAdB06cbANpC1gkeyuXGXS9kvYZqDG5HdoNpSneaoFScddkAnXc+OX
TSZLrW/l3pNdQdxnHYAQnzrSfj/RPM82buqzqmKl2LdRYX+xZWloMZr9TiDe4vDU
kO/kUWZOuDsik//VKsRZbz/zb3+v4yViTSCztYFjcfm+VJX3WjfaGGRm8u9tbwvo
g8wpH9V9asTG/2nKAvvWLX9kMGQgfeebsALwrVWw4pe8NUqRRFVTvgpgFIemanhF
yPYN8gVGMJDR8y/QlKfcVTmvoqNoCoe9GZI3IQ48lQBzLyM36PF118XMK1OsBnTP
nokPAEki133BEGeE/RkFmL4njDqvW43iwCGzRw4YsALDABqP1zy+v2LMcc43vygr
IyOqoVr84hxVEmFA8Kk8WmfwlMB6kW1M+g9s0+iAisdUh9wAJQr4lujGRXmo/EwQ
Nwz20jKuMhK6wp9KykrQlmWQzAnppeRit3h7aj0FXTB0nX0kLGXFO/LPvlC9QQ9y
d4C9g9czNBb8qerrAOzOoFXnF+IhoWdcUeoOY1aFKi5zSbuLaisS1UkXQBOpBoBF
qlEBGjUw5rsZBAk0Pkjkav9uPI4uhOCVAnNw+WweB+IgD3LqkKHtYk03wGvo8CUS
02I0Af0+yBtU9Dbs38WhXk2kNo0ge92IJR54FAxMB8UsTlHaWuC011X2LR0729P2
1Qh6I1Bb/kBOdah4FvTbEljxHv2NqGEN8u2p3oR3Q/RCfflK9WrvXIWCd2ui2n2Y
5yfXTkcKgh3/shO15ZfXR1yKzstVxudmv1VEWlRhg+O7zDaL4NX9jwq1LDZmuzXF
eUHfiIAX3Nduq2FIea9B+6Wo2uZEVIf3Sjgl6Kga2OujfSjSRKJMdzMT36Etglz1
B+XvZhru/liceg4foblaSu+J2LCCQ6mlcGPYQFk2syzXzoQ4+WVSZ71w04rLIYLS
uCzs56B2tk633iF6wn6/QTyQqw1oGerQ5BV9co/2x+48KEYg0FQEi5PcV4nPtXC1
MzFnUm8KmTQBrEliBMVlJ1a+ANzt23ssci0B3z87jctQkyHtZKeY3QLLUG9BUEyO
qIaK3383pVvkr6A+AJYqO12LFRRluWcB+juv/1fJJcSSt3O+x4fc83/6ugA6nHVt
jxpfQTy9aSGZXecsfpv+0w6kJ5HrdTa1MsrGYQbjqEgkTGQrSPBnt9yNjITum3ep
KN51B1W1OYp/hH0Em9BdZy4dVlH/TQDLZUhz54CSgn/xhxx4qff6L1fE4Gz5jrad
bgt7XdBWX3eXd/FucCm3NtOIl5FvgPAKVl/7ISwraFlQKiQGcrNQDHEky2FbkqqF
dzx5Triq1VqiDwwl3axnnnhIxX8Sg0SG7KD9V/n9/2x5f6GhKEC7NZqR50XNmSzm
loIWXxNTShI2vHLYFh1Tr4ptS+gLp+pEIuRa7Gpr8RZQAUaO45oYT2HSqYU2kxlE
6CMVPg+COJkQtqXDZQMYnBU/k9+dHsSlKsS6S4eyzjFY3g8dDoG9oUsi9Gh77fzn
qqcNSOdEJ1vUO6JKOj5lumGUZJilNAXt9XmR+Ean1YvsMwr90koJ5ALX9mnEqIce
DzYqIdZ1yCiaCs4zPEWJQ2JtPLsi5UNtBYKuwHHHKmde280q1LEpTVBHarikT6z0
QoVH9LS8d1Y0xRcNyIR42OZR7eO+OFQyLPH2ITDG1hYttmKrzEnEhv3syx5PKIql
PZzPjErghMgXQ4+7vK58m9OLN+Fi/doBFgENArAT63WxFm5aC19DDS/V2A/cBbEq
s8kQfGww0cHryNp4ofb54qcyhocoEh7nWYZXIE8ZIT/wJsNg/ZRw8wyr1ZHAjK6S
wLH9ySneFdL+1bkVOWKdZuCfwdebRn27gfgl8ZNkTJExhPsPn4r9WIqfqDKV11ZK
wT0QObsZBz43PrVl4l8d67kvI///YF4DxrCSWd3l/t0YJLwxUPfuD0uBTHv6bRNt
ttWdX4X2xOp+Now6EzUMCAnpXlhacIShrZWecnJ64ZnDQXPI2hzLx0T+PqgHZ9UC
TDHipWs76eV6nMxr7OZ91KGL6oDzuFDOP80G7KTGdmHCOp6GmblSPPyVWwXsVUv6
Aj2JwHKmvKEHL/UDW9nSscX1/i26j3WJ8T8w6Qbwd+3ci94c32V6HKDSPWcnZSEp
zjCrIBI704DTMOTj+vm0H4lyRo74C+MdVt+O5vRQP1ri3HKu7muwv6OJrzVxRjWz
JPC8T+ph2oHGMjVUa6p85U5KFuBj9UkIcJgP6XuVVca1tL2XOO3eCbXMNOvQj9P7
VvKD8STbYqnAoljHftakxEkUVIJ6A7w8zKwqu04EjjyUiF4iJ3EQtLM52E/Ug4WC
y5zD/zv23+PpAqNUlaVaigHSiS21yQRmvjH0AbvpSG6bpowbHToE1uM4ZQaTcZR/
QqOpZn81/0Abq/Gi2o0kAUhMBIO9ysJ23VlfahUctd8BEAdHh07rcqLf7qYPEVHg
CS9JKFk2C2R8waaBCO+wbW6wMj8nBrvCro8Wmog60OD+WSRgUbZbJkBydsi+f3dM
EbUuX+uVniKElxRVPQ8RlNmFG2FU1rpXrigYVk2L2FxYftJzvnbFqxIlI6HdRj0m
o+xMW6N2FC58ErKON/BUZU5gpSTtQLT5+1ufn6zjKNdEXKLJ0uo06yuR0IKXtnpp
TCVk+cqqVDo68X2RrHD8+3P2ZPc76ei6nEpAmLHpM0F358PFQWsBHONGCDdxDZ48
LaeVdtUaE+thLoEk35WTFOhZAE6VCQXOM5eEmiAnt8dyGcKs2EmiDOKzN3Kohm1E
w8DFb8LeZ4att8nRYRqsn3O8JxM+1Ken24te0VPCkIcnHW2RGHIvl9cN6PhhCzGs
i/kgzr8JfWBG8slN6M+eFHEXfXWD9enp6TRHG+d6rHGdVTABTaE7GNy6bSd12fsK
L5EIHpP4MMBnrGmRh33mymUJtzQBwFJ8yV3LbxYnk+d/1mVQysPL5ICMsure+vPB
Yc7nzcQlzFBk4z+eodeoTYyxP63DiU/BV4DQtVceAzyIi/xEuuCCvOry9E3aeivR
qfTFtLl4TEND8dkolAh0nBBXfnZJ4VJOwIURImGasAvtxZLT0hQ6KJA3T35CNoDa
HmLHBpu69F0arWj91oQLpd1f9IMQRuelAoFnIy+hQCuSioozqAFPCTBc6Q+EtPct
BpemVo05YCMnc0eV48tN/hf2Mj6V4qKRmtdNWVqbGg6N723O9SKiobK6sLYtAYXh
wMVuXw7by6C+A4YBw5KXfmOIJwj2vEO8DQokbKGI2SQPPIcjxpL1C8Wf4jtkHG00
jVw9qp0I+3rwSdika9OVaFnvF4JQOGCVL8X8/MpvUi23/SFGP7DQ8NkklMhhjcl+
4+ubAMSu7sLMO3q97pqnJvC2dcGifJXwv7OCWu7jEShSzGGHmIPX2olLG8UlL2Y4
VvlPlxWBScWyildiq8k3AaLeSjNKwuiluYRqMfMMzt9ts71ZQf+zH8pQ2TlSYgbI
sC1mtF1SUZt5a9u8e8ZA8Q5dWquGFp8NarynrVThmCFIk3ZondXarW1YqdTxRFNd
jdvXgeotbydtLb7U4RDutCBavsD6Freyv+fESupvCOLR88nUV3ddqOWjkuQSdWXP
Y9JxhE2xFW/bOl+Y4iquIJfygfG3PKDMnEQvco9UmKCHfHiwKeCPKnNDqSXTsRfk
a2epzTJXcGBYy9uTnsTYR1pUa1gIZq896m1NR4pyU/1W0LmsiJVdq/0UEfhA8aRN
ULY5gYlmOHHMu7IsPe6Oclc1wBDT/NFpSeLHfePRkPAL0YBU3pbIb+4/QRxA1xJ2
kiYE684ziHYgC7WtKLoTTtqpJDqsMpiTxtf6F5cBSID5ylPOeWdzq7qRp6BEKzsn
15rgkRW1s/YfXGFHBX4/UW9ojtt2S3bHau5ZlIKjZFZseEx9xv1NswJQKRg3H4Y4
bnsvCtDM+Yiieb9WiDSzvxUSJtJyfiZIKPHMuga9rIt3dn+wRLXW1UHjDJnCDsTk
HPQZJI9GP1yT5iklAnWtuxJEXZRz5ksq8VZ0SuxZotxF6fJbJNWYRzf43XMMjoef
vrFymL+Xz1Ya98+n08Byq5LackFPGWkH1HwxrCRX8ziPEUO66fBQnW2OTD/1SI/x
ag18fEHYaA5x769vdXHejBMYHsf+GdSCbxzBxcT7328yRJdERRR609T+2sOW7dzW
f6nbmDq8JEMNW5nPjP0mfoOuJPkjqT2FvrW1W4yBFiV2t6Mz4vrsUBzRnFk78xrj
o5zo5zjaY3Xa4bcUMWZqJevSWT6JaJ2pXgfiIi23AIjHpQptcoB9jrhs4QIJ4UGi
3tXRkl5Ipi+sq9p4YEoL6xipCUUz6o5ZOnKRws0NmwVddNdqDDp92KACqjS5c1SJ
5s90meKXQHXuoHl3pGW/TdWy+Srdb0DKVsxkUrBVWY+xcHIf7ijmkynf3i5eX9Qt
RCFuRgRUaZoob9J7wxydZ0dpQm8iqQyFh0mZrg2KZI/mchJEqPqWDEh2ms6NWmhu
JldqMD4ieXXi5Yb4tHGzrKtsTFgklRO26S4EnCKEcq2tRjsWFO4loa+0oFU+oEp6
9kVoawuHb8m32ieSu/37w+u0vMpmJ+gRh90aQEmX7wi1veUUM4YEpgZpuBBf7Ytn
QNnLnl23l5MOddSqQR6hyMZN9en6n82au5t8hqiBo85XlFavR/E6qH9CMY6A7zTg
4U/X/AacIq9bM5TZqttQv8d6uMd/gkCImh1dwR6CCpBEp03Vi98J49+Q6uOC+nZB
HpbvVa6Gd1BXYYK1540x0k5xN6mLQ+wkh8zDYLL5eo7WVMTIGqxfO1PuKxU1dm21
xK89iDIOse5TZaxmN3GcBrH7Hout1WIHkz3vfzLg1VUNqzF5kcFVnSbF09kdR1zp
kE4yrgOpv0dVi09dwDTpOnGrWqIzhZ9aC5aozJW+KAHzQcSi6modgeXgp1ke8YWb
1EGiHx712OGWTwBlMBqTk+vmq4FK65qndR2OHHP/f58cJMRz7AfKL4CzJ+XaiJ9Z
fB3Q9gB7OVggMpLziziJCTdsAIcECLHJmbEoz3cid2eEBTsiTA5rlfkg/ZiH8HRz
OiyclmZ4jEF6FrzBBY2wOsP4v2H+spVGQzMl+rpE1D48isf8ByQqGow8WX6ul+SN
bbZbZ8zUqNoxk1Xn7HHbsbp6Z7bhtZ0R81SKS49edmIgTPs5AecU66iaWEm8vlz+
ZguP+B+FEz74f0e4IstdUEOvd+0olCQm/tx33BRb6zyR+1UMqifHHvNhOpeZcVrA
oXEq3dzEoP4emllGoEQh0ADCry1DyA9+qd2boi0H0GysFEjrPD4A5dib7rnjqyHk
xB/qoE5ZZAaFpXqyi2YlTqokXl6Wv0UBChhqOzBjueblF5sNa7UE3eQq8N4vnKF3
qSIh6p2oP9lNpdopfru9BowgsQb0XffSQWuyMfwuSEbwV5J+KmUg6Bf+hnz6hAlu
tE8JP5Cu7mLkrtIt6VG4b1Xt7q+PLwDa9TQGluZKmvSRzyY1+jiTrp6YwdGKKMpI
bFmhsA+V7G2t1gN7/Ag9VwoIGJkZ1RZDpG0vBkdA0xGL9iA0ZA0azz3ZzZeDZEhZ
G0WU++70i7LjIkgxRNNWjs0579q2fc8DA9iRjS8M1BuiM/CwH4sScqX6yyh7ObLN
kIanomFHHBCkO/BWdfVtp2/MIluIZ3WsAxBUUSs4RFCJs7O92UKgq3K/oM0Zs6v0
7aZkuqG3qVu/7YgcdTD+DpXE7vxBflPpVke7Foo7aC4dvrHDcwQA/r8zkmKBab1Q
X1wR8xKrlgknW7nlZI/hNa7ZyjUIPmNWlc/VHWUzftQ//AlrtlzkjngaMpX/Zwzc
0fJnvufxolQ41A6STZBIohcYjHRRRjCzLiL2NT5AYOXLnzMJQ8gItJhPB7KSXo5b
wJVre8/vh/von344SEP/sXFQQe/g1WkOqAQsYqc3wLlr2ivIr2puie8fW4aALfaF
wc1HCsaEPvbqM+NtUdjDEuW5mZ+fcR3RfDOd9T/FrFkTKBPgQ6NHZnpFyDXGXMy/
SBxyMVex/yUdRYovnLSVhfNNEtimvhgqQ/o0XE3M1w/M0CJgw7Tr+2Z7ONNhdSAb
y5utrrnHOQBdhw71w7O31M/BgXbTIghQ8nhyP7yIyu5Akqw+9XGB35zDil1yUsrY
K6X7VRwD6MsY3Fd7+CvAEFiyzKDyLjEyIFLmRCUwC3wSjCQjadrQEI167igE0YMa
ECqZqPL1DKmOqHUp3tjVhWT4Li2TrmLJ1jRNh+QuK6NE1FwTThPP0ZrQ0QoNkLje
1/J5yEhIJDbbqyHGGH1ffYI2rPuMaKjSa8dThQTBjBJ9/jXc1ehZSiBFA3eRpDnX
bnqfwpfHkaE+RYYQvU0uw4BK6Wpqf6ky1TSNdwIoK8cbVhp3k3NU0PJ9l7WP37bv
VUUZm7UfuFEcfIREWNw3v0nYlnOlGAJAwLyGIoB6j+UgzN2ZA4c9iUvS75woWx/K
I0pFGSH/PiwW+Ru3cjItItu848GsDSSMwGqxXv47eLOwW+0xhy9fWILgyS8VWnSs
bzqUj6ZyqiIAQAt3cN9M1HPLe0lriuj0gusUQAtTWmZUIjKeH9vZuQyjIYir9HBU
usykfo/HWnehWBmfWLMfzuodfjgdXtkNYAyYmllV7VthiVJk6TiZAFayWhgYwW4S
Sjl1knwO70umYdlku4fVGe8mrJePrHBEogExmALR7b2dr7W6nwBsyAgfnAbylYZr
kZgcI3AkwOISaAA79D4v9zRdW7TATSrqlb3sHiCutkh+eovexjZ2oZEAHEP51IID
RLtJaL3ckB39dCREtqaaOwiRJnbhv84fi2txpHs7j1SdNu25WrfOF/2i3zv5EkyP
Tf1wZHsqu3egzDE7m3xRExuYqaU8osNe/l1gw+GwSq450dAHWp1zxGGKJc98jg1Y
7DZr9YLD9be+R5blA3YHKVKP5j2r6bYoRSliwBHwDdEjb2Sh7qlV+fv2cNCRxFfd
6CmITG0dKQ/+37YJIfQN45HWE4WCjOU82aaWMxzW8kkQvliJeNuAyqPj763ey5Ok
t4i5sr9xgE4uBd8ibAbNqT3pJ41BcpF09MJ3MFvPO9z76+z9lDph6xzpOmlmSroY
m08zRnkxbjKHq1nYa87wEiEtidb5wrbcXffPlr+rNpGRldgxjQw7XNW+qqyuZhwH
2IXRJ4YFQ1/0/nunt1TnCLF8SbPNd5vlpwiBNQAM6hkSkqekY6Eykz+Ab+RqAFbj
knkHYraiMSbdAvm4nmxOp3zNr/tkCfedRn4yc292aQ29+DzeoTGAys4HIEWtawgD
swSHGLWZYWGefQuwa4HddnmTk9g6u0vSw9dYqnagYNr4M8jH9apAqnPOSYhCEq2b
k5HRU/6bYBRCGpPhFX222JTXtm0noJ8BNodIiW5aJaY8KXdp18cShyVGn7IQ+g6B
waNtwlLJpWyN68Tl/8bzlaJb8Dv8dPwLGzBWl7HfKh7UIiElSZKSra5mzPAgEvPS
6lNhSXnX5M2iv5XzWfOklKy0xTjFuEeaaoevJVWg14pXSmrH6zNGsnoCQdk89oqj
iC6+z2h1SwjBzhf5VFt8UfDry4XF//gFZLO2vtydZ5LB4kS2P/Q3iFhVnsh0cTVe
5y1Rfrxi275ONoL2qe3hNlU6lnIeblV955brt6IfSCnvcvBusc0E8CCk1+FHRACp
yXx7V+90de/9qHlj99tl45h8bi8eTKbaXdS7tl5MveiXR/tB8bnb9P2bCmvtyxW3
saGfsJyGPaIW8CpO6ih9bg4Sp5/DkkugXLHvWkwbdCmwgTm6AhcS5IakxS/BLDwz
4UT+yUjPGOji4c3TOeSb+22sbpTYOu8kD1VMi5V4+qFGafHqHjVtd4oezfBCOfHs
Y3Z76ypfo8BJYZDkEVNziAfTFDBOnetzD4txokvYIzjZE79ixMuBkRIrV1qZvwy2
Uq+0G95ikrxUvr6ywMBUC8UgLNI45Gln2sIx0YW2eKBKK+H8XYeO49UJ8+nwK7NB
XBsCKxxFNsZenBuHOkP1Q/sCu0DgJTK7e2B6e+im7Gvy+69wVz4EXrXcKaLrIjuE
vsZ1LWCNcRqtlu6ns5vKafdyLG2bqt1fv2L2D5+mnS9mXHfV97PC0FmMySjbHpTp
n8xu2iFXmmNTuMq+EkTmcUEVCQB5OYdX9moWtJFq3iHk+4cfQ6RwtiGqWAzNTVs3
7fBjRumvo7mrpa8+m302HFO/5g8l1+31p8rtW9Tbt2LL3vi1H92L3OCFMm8dIy3L
s6WOs7KOJ/jQr+1p6Mi/BBS1PuZgbdqtlpfqZBFlF0GUvOx5Q2kqzgOwrYGSY6Ss
iFJ69cIDONWDEhSUcURIxwdfRwX59DW/hdKeKwKT2b0IvH8b+ONf9MhkNHKx5Kfa
LbKs6l71JaPM+l0AMxoZOEhmynURi710pa37OcudA1PQ5+J6nJA+5AnpCY0UGq72
xkdsQHQ6O9uyOikzkJuDM3sidFgKwkPOXqjBI/kWdEXjK2zLnM9n/Cusxklv7rNL
3MO7X57cBGJZPzuQuoTUJRjrE7f2IG4TorThWu6N+XhfmstMiCgPYgTxaq+UiIoX
8lHHTsGoCdg1mW2jBJNT0L42hPmslEfqXFBFLZ5RPDIWRbsifBhj/TqdPxaau82+
kg5I+1MXblDdBFqPB9qUw+KOhh+qypv7OUXZVpkR3fsl1CnKcOqoimYODhiBGy3t
kDXJs89MoRmpHuh56wxfeiC5nhIewpyCRtyigTizJLj5qmR6YlN/ERPPPNF4GK2u
x0lx5UYPyhLyqkFcaRWMi85xOlmvP/4nNUuYeAYpMPr4diVpBfrUUDE0ZEc05sOH
+8DpQgC6hCJsZflzsRyGO2d9fIkR85Wgat8hqpLajhHQecDtcyxzanN2AoD+rz8O
K/hcT0/K//uTcXp0dIxvuOs8V8Tmim/TFhh3VlvWTFey2hc5+YTiZO/nkfpWEvUs
FUJFBIjkPn9ma83yhGQBsgBgoA7Gv3Wh1pShuXPSM0CfsECMYeud1SNXe9dLiD+j
5213qYYmWK7EQ6Tj7PYmUzwG/OAzAoURo7M/qCWqbTSzdpg39jf16xjYZsP7I51E
sHpxj/x33ZJuAVdogW3z2EhKz8yYMF9e8RlcFjEXCOYPetyV38Sx4XPNGmwIeQ+1
4IwJjc27LXf/DJkVgOSKq7v1QwU8+cnAEoKW9R2Uruwbnu+TOXHfG9wsm4QsDPjC
WOvgmnlzVdDmiSu/u9aRDN+q88Bpg77Mmu/n438/0wwW9Hm2L0iGpYnlmV6vwR9Q
P5MUm4P7QC0hlRa1DjqVGFBjtiT3qP42Dhim9924tppZoG0ZpCVWD7xiOTBA839G
4JbHE92FjOQ3kZAgBUNnllxUXz8ZoobXQmEEBV7hL6VM50uVgr3y6ygn0gXMfs3g
ZgZYzlV9kkuKR/Mvqt3rLh+/0BIoR3lyfCndCv9zC3uQWSNhI6H0Gd84TZEzRf4S
eGX55eGMcTr8hMWwRgA4OEuTmA9C/rgLKv5JGNaJEijpwpIY/JrzpUaixRvlVuOU
0Du7VhdKbkra+7n98lc74t90NMo3ZD6KMjF0yJ1ES7pTy20kLwOIejNTtgfDioEa
vRS6iXAbbG2SYUU0IW96rXGaLz4vaqEbMUyBHvq4nOkcKmStam74WhY/ih54BnwJ
CI6JltQFOEFz/ONFx+ZqnrrpZZ0tJA9kRNQ79zjmD7ygDI+dw3Pm1zsrxIGMZja1
pFe/929TOAH8JB9CHH3O6+Lz/MVwUNm79h/dZtaMd8V7sIsGT1gL8ZTSxeAmR+f3
421W/dpMOXc2fhRQwBRxxnkE2GtD0cHe5ty1KPqDrPmSX3Ugm0CiD7bFaTe68g7i
c/RQJ43CeLjlA10qbDbrTQ195y0nA5n776hT5+fHVeCiS0wVh1Cv76NmvW24dWRb
vAcwaCxEezrCFqVyxqTRwCi9hV1OPBzW2+85oGv8i6u3fH/jAQvA0yWBsRCtHJ3M
r1ckAN63BZVFVuD8y8P3kI8SMZqJOmkYOLOKQFXbkt+SZ9zk4ai/WUVx2nA+W47/
ZqqdgoN78jxAaa/1jI2dSEhEjhMpzh8rtb114EsvMfDaPfSCcLC54lPSgcBb9cYV
jvvVtjHNeYZi/xyK5nkMlkUT4DyxgyxqmnBy70rSJH3Yv++nvGGdrywAn/EWedvJ
I1PeJeTjOyHRUUIZNNU7skiuap7EDiGVyGqLplC9GN8jSzu0tgs0fj9tQlwNsaVk
uIc3s/kzPQWVdp0PpC03sTxPWnfPb6Pa8S38YPzg04Zas9Ww2JEderfJQc7QNOre
dkyP68JtNtqTFwImf3ofJ5RbVDk02yiNiy/yLbjF7DRMbKG0uDojYPW/vHzBLYlp
PPGiTYbXbXctlH3pc5jJPNkAG0wgSwRnAXptu95dZjRqVQx84JZBbTTQ89QLXr2y
3pUhXMMv4Pvh6tJQdhuGh5c9ZKVrT252IIU91mNCBBmkr/NQMIZ+RCvq6JGSSXU7
+ko64hNAzXYYNGdSdl+aO+TKUEpoXLl0ixWx0ca+AYZHpqVXmYbMPM3ZRnZayVVK
C5NJfye45uGRolxT600OspLwvpvvmEn374MjCVTJBOxAmIqQ587mScYtO2825ZuT
ozT+/rCNND8vLdnseO9qPIdOj7blhqoVdmdsIjnkz4C0FISf+WDIPtasxJyGTwaP
r1lbPAVghOTim4QcwgrkIadDkNzKDVzEaVziSaqlWOATK9oRd1rWy5q3uJ3xCgdQ
YoKlItaUv7fSHPxVw6TYgKM9R5cDGSEG6lsQobS523f08q3HirSaoPdS9isfZ5jG
eYTFsNQJQafckV8BHMVoMV+x6963uaej3BapePvqoRjr0IBY4VPeHW8T0qoGpZvG
M6rbfoG6qpRsVyf4JH1N+XQ2mAF0FN5zi5d280Eb3oa2Yoi6p/QKsFWueVDuYkLl
PIE+YwsnxOkpfxeBS6O4WsLBiEqXeJI/Nm7/PHJIKuGFGqqoWJ/b2uN99xdNKPpS
aDcKVuH6nkdDCFh/wNPKHgZsiozLJZ732HIngCYV0QKx0LLm+oMcjeoC+T+JMnL4
NwDIkzARabpGsfFSGUv1U7l6xbdTWSuA8YaB40x5Y4Pn3xYqHcNs5VSfYcy4/BrW
xFChK3kin6ULaAhRo3NA2ieOqZDvQw9jKLABcc5wRUdPUB4fPHXiJ4CEiw1k/Fcn
EA+Bble3Rv6ni5a1YrMChT+OU5RsY81sZ/+2yQgU/JvMMyQjfBdcoH//eUxCPiY4
Qe8i2uNnLOnLMFay1dkzEqPuJImQbgu7Mwh6ZHN/YC4NzltaUdJANkOx7f6d0ezZ
Mn/7tzM5m5RSCDix0eOA2qKk84c/QeFJY0CXuw6pj/ZyUdE/rRM8ake/OLWWUF1/
/JyJGimAoirwOgh1RUyyGbwUE7hIvboj5nwuaVCn9qGMPl6536HR+Him933t2zN6
S2saJONJhUZyaSaGlQAhzigMqDcC+d35DG5xPG6kJC+LNRMnQv0St2mAV5JcCzjh
d3RwpCtHnCspDytYsGdPQlRuBWmo4n25/eu6+26vZS96h2FIJLzNVXUI1wjLb9W/
CUgB1yTZpQc8+SzjdsgPnyTTFn8eSAsLueT/sIaoTObkASC8LY+Bq8wAQ5qlOh+M
5yD5uZjo5lxnumIC2hsd7L0NbcZ/n9oLxtfI0BpU8/T3ZU7kMnsi2oLfVWQv+iYA
NUYPgopYxpldXWwRrKr5pWtSJyxZDrdBhJyAylTt5tJ3MzRMElx6RkcDN7/n11P5
n3RGDnjnvMijJXI8MWhXcUSDYQQGFSVOOpPV4yvjXm5vcRK5+USS05bIMFiMhsdG
K9HntJeG847is7eSY2vthPwLItS2h3bel1BCL/SC3+C02ngc0fQFnaZ0PB9jcoum
xN6gDGYbSPJoLCfwJRIXI1RKWgZp+nEz4cKC1uLH+pq6fxuim3s5fmPPtlMaAk94
mYxVRYboGFJpQWVsF6WFJLkVzMSOWtb6F0aZL4hZtxRbAy24Dk9/stvhO5FGsNGW
IZdhU4Jhrqwlse99oCMlqtnh47sklR5KDHuHNqMjZeYGhAACJMmx3UYrmoJCPVk1
/A/Yz5EP5dueHHeuDaiKHsFHA441A11QowfSzSBpcq/d8KDaXwb+NjIGuVd5Ntnw
glXLXpL1KWvW+ROox/cdg1krcwWqAasHodYfIS+cnp0j7wAdfcMNimOsQ5pNScLC
zmXTJ1psqj/yrbCgPPi3XclCxJ+PuToyHZqOdxCW/66lTEqqhtTiy1Hy9Yd7nbnu
WssammgYNjAbZAaLiWfqDe5ZNtb3bcwSvTLW/XbC6beDqjY5o5GXGBfxvo5kNGeX
QSB2ye2v5kbbDxP602hVeDr4oUntufrM2fRQw3nxdxbkduwy1Re56uNEBKCBYLa0
5/0VJA9hvTPGJlRmfErNRgdwMogoKiUlAF1Fyfo7Q4dEfpfYdIUNIZyn4odA8CWH
YNW8RbiVN4yBi89Hi3j0gDdVI1+ByupXrHUxEfTlb61d8guOuutI+mFan6BkaPhZ
gmjKx8s7eQxXfdLRLLcg1BNDyoBSN6UHidf6fSAh/fGORxEHHYoWqrbhoBNJJepk
KfmeJZZnpYxXF54d9ZIn07lE6ks5rY8vioBrbyufk8rb4kLGatmg+MmKsJJ3xWkA
/+Yfd+SusQrRohUmVJm/gZEy/h3RXwTqsTVJI+nMytsn7A8lP0RwN8GDVAg0BVCH
C687FVmgdgjbYdGFQdeTyuMLtjNX84HeQg4KhlYgC7pu/Ck9VLbKslYspk/ePbp7
/zZHmEl8hQRyCMPjy4cLWF9fIMaWu1MR8fmUbdC4wBmfxXuq7wZHpQxX9hI9tI7A
9cKpqxJqxyXPZLqW6pMJ+tj4wz3hOUOEdGb4Jr6r86do4k3/M8F2gXuDOCdKG1Um
DqTBPwwln53wWRiL7QP5tDnYZCogcoIQUf4DA4azgwxxe9vVC5SoxhsfCz9NUD7a
yWrEl+cJBuDNUw6h8+pey1O1HQDkKu8IwriOPHBHJ673aAq5ijWnvKRKPIgyp0jk
Siyz+9FkSprxM4REokeJlaGPshzN0LqJX8JDBJtfvzZYPBBeMXfuX3xf89RlWWUo
ueBgyydAeDwUFjC979N/RNx5dO9GUb5rdxPujSsc0xknoQlTRc60hQOuQzP0mwfZ
KwU3siowHB7ikRbTGo9v8K07qunVdvZQkaVEAbnLuOOZgDQmi722qHkMsjG680xQ
5cIS09GMOfiPQT0o/TgWpWOnd57EZuAKctcRbPxQU8g3ehnR3Ewxeg1rJc+6HJe8
ycZ/E/3oi8rHoA7pZJY/Xd4IwtBg/tX+e7jH8VKJmITdw2C+XcYs7ndDJW5dc2Kr
1yOVzRocVx53E5cuLwjWufdzMhLyYmSflkXuGGAYpvsZD8XOxrX9S64b9BIA4vSf
/hwfrLWNEHcKZrFUifZ44926QG4/oXYt4k/CEcEjcFJpv29n6G+qvwn6ZA7LJfpG
DncX0Kou/6c9Fe3k2oZXaL0CVguNkZ1lpwJpM8LonpAYIcD5jiLueMzQdLIqkLTL
xyNU0kAJjYVTMpqtafHe8+sgEKkPqK9QAyvXispkAXoH4gZqS8dYMnG1Q1kmvRMf
cz9n0lVZuJ2G2YtGups0HUw7o4ozYj6CsAeaDppDjaEEoEbmoi62HTVkSf4sMq9H
a7XJ0gxWnWt0SZLJyjZYNbOU9oMOHrtHDWIeR/ZDapVUZ5s8voRGe/vrWcucJicj
w7TFPwafSD5jSD/7Aoen3XuGyIs2AGI9jNU6bI1y9M+Ns9uL4Aano6pfUMAbxWKk
eAqvOL2rLeqUhAVFMV9NXz/HniMDloYjIPqnIvj5jTSrFsS/jKeptpJJ7z8u7OWL
33zYt1DrMF4UxbThXqXkuKk5oAHryurHRptZ66Jx0dlKqKutYVG/QOSgO/nnPYQR
6rFj/2D4sLrwxdjI9oR5ECy3pUUvFU7Wp/OPHttd4Sg+UggS5liUpcqsY0YHkvQs
SiZzAoZmC3YSfUYSW4KbhEgKcCZIZ0TXjo7XyLUy8imo0I85gKZ8dpNJHKPfJAch
X/OvX2YGZUaYSvvq1PI9kv8kQSQWn3UeVBHOXCDZ7VjS6IJnkVfJoVzB6oMyDQM2
XGQI95sJq5Wu88in0OCma6/PJ6sVrgM6pnZuJtzWzt65maPQR6cwiMCoUyUn5Zez
WfOMLKLeP0C8Lct0FFk98r+vsgMpwo32afFB9jFDreXIiSBHgk0ddlLYQOUcN7LZ
4t11AxihCja1NKiZy9HCCvzmwAZFk9c0b9JXv/Kxquqa/zlP5f3lHRjv22msCY/D
xJ0WFN6WXlNp1sbCPhpuMJ6YWZciRZ/JZYa3qWU0KFwYWlaEy7bFf3MNGxtP9/wk
EJxLMPGiP3QbGGzBguUQ4r1jAQTiZL338ECsf3nVH8PFfnKwfseaXzd57KzY677x
hQUfuNLGkZ3bl7/4V0h+lhRtmE0TzuiVeDb8t8XNPsqYK7pF0RPkU+v7ZazHr5IH
Eo5gUgTiXinzvns3FL2NTmZshKp75SqVwLxUsUAGPk8Sa6dn+tPDJD3+oahdQcgZ
E1eImY2yHtC67fFHalpIMBzg3BoB8AFL1POLca2U6zIEuO9k/azK4yqUp34fJxJh
UA+V9v9ZHvqTGZKfCUHfp2JPIz/gihIOOYaH4zCuf2X/tt7Ev+w5jSQqhgLABHgl
o6XDOlV/0T3aAlq14jgvBDENu+AyMZ6bd0edv4GPx6VO1JFCXEsHUSVEe+oct6qd
6pjco160lDuIAqmaN64DhZ/NCeFJexunXXTJ+0HFo/jFSQGf8/BzFZi5is7jSVr1
rkkfgy3QhxltREXdJGdE1xsvoPlJ6NjpFRCr03hZFm8qBekkiW3rKhIY65VSIbaw
xX3NODrTd3NhSBDlYK9/juFxeJhUChlZcBD9lLVbwqSToAUxCe/vNpNTYc3wptDd
XQAHRzRdICkdGc0YKcZqge8waUXVE3JLgHJYcReQLOn2fVDF7FouYUbTPfzpryYN
BSDchl3VBhgVCQyZColxVHd6JIXte9Lpil3i3Uv3217qF1Xxc25GdDD25Pyvs3Wt
oRtr8RVjOa+K6qZSE+GHRKuIa2ZeIAgyIG8VrbFUI+QV9x+8UxAGG1wA5splwc2Q
ZtpZfgszZCHKDMPheH7kKHhVbb07UV68CVRLBQnmfsB1YIurbzlSiIU0LXj6G2YL
LqOxhRDHl9pCw72sCjod7j37+xVBUS/TDR8M4LMCqCmSfOQ1qE9LTsabNN0WXT3c
/wFcPn5b8S3z2EdmtiDQIEjTb9hyWSgBmy8octMyYdyq5jW0fUC8F6TYyR18BqU2
JOOlJ6pxU4SXULPR4+bpKqrb6eeQRVrSnMLX/5UmVh5Ng7SnZpGQpk5l7VCTDpgI
GT+tlrdwDEm9O6LjZRnxXi712x6tUtQSLOFqqfFQa3deBCYBioSMgLHPMV5bL2oJ
LZXMEcblDOupKqYYm6pAYIQ1l9AaolLFjsS/ro126VwMXd2jYGVP+ZX9WMlxao3q
9H5A6OYeJGEVCQWLY3+tQOzt8gXGbxq5IJ/df5eg3OT+SL81NzRYWdi0ecpRnknD
QNcwoO1vwHYfbAT6hF3HLNJnglo7dqomNw/RoYq6pHZ2VxxscPpocY1clJde0lCM
dDUwkD6ckQZYaobia5j+XByWpF3GgGvuMVzWfZehAemxSOH0rKWgUqQsAeCs3tDa
hmbeVObU6bruQaMiH+BaGra+/BI2b6wQUHoV297hMm1ZmPqH7E488Qq0Ja1vpXDU
l1IJz+dQHjj+enxk9bPR9H7ncTg2WTMSqscBrTnzO6Qn6MIp4pFIQDVgYuckaNlK
z8FcMo1AFcpYB97gBkhVOFxyW8yHyOM8ZrMh05MK11Bjph/KFqsKr23TwLvC+kFC
y9DYwoPUOPDNZKoyuYGd0betfJkKtpxFvlRPRVDOGez4dVD33/qU57T21Zm9faxO
0tXRnxCgGkE+VaHERt3oQ4vYen4ZiK1vP7SIYnshAQzfZworNzBsZ/ekBp9ZlPyK
/FuzHCUAvl0q41WTkPjkjm8l/cFd6lenazZdXslE74F3mVzdWU93HYCgOguGZH9D
5Vhrud4oYNc5nMjvyGoTIBz4nHBq0xWSFbfx2EvGsOQBIfxIhMEkzTIVRmHjDW2u
NggX2DUBCp6DLjGpMIlTWxFV1sVA1bYMNt4hpztuICQij1kifBzwWpDmHcwv2uW6
rHZT1H3Ucb1JDtmqCEgwasD2SI+eNHfFIYruE4Yod9OoNWtKKkVrumNnR/pgtypL
rrhIu5uSrKNFDwfpbEbA5sWAGxjECwSiztaRT5u3YEe7KjksFh59Rsnc7AiMVvhU
XAVC9dIRZ/OPE0TjnNZnwQEpZ2BiB5uYFoAcdYYKCmslN13XFE1v33WB1+AcFNce
Q4Gn2WdLJssKhuuRwQQG7ap4E8BDa2qaHHjJkFLUHxF99WVjCHE1DgJ/dnL176sm
9b0A10CLp9CEbUXDiZVAxYO6UfOQ3WyO+fwFTi8PXO930fSwWtVCXeeKQpz2aDPK
1QSZstSDXYJMmzDWdAX1PIyEIYY4Lcw49OgcHNlqZNIZ6IdrA+l/lQBxh/DU/GJ9
ZI/h9+LaC8IqmgJ3H1FqcwRPmQ6nUj6n8Q54wgQZbIhkF1Th94k4yqJ3yY3TQgYw
UGNMVOcwey6V4XIWV44/tda/1+b5wgO7PE8ctw9xCjnJRSoWha9PbywGKaOIL6fM
ilede/c7hX0q4zuwLWs8xaKYgxLVnudXu+oQW+VhM+VvklJ3i8cz0woHQXEy+DyG
LKB5BwiPY16/k1vbrFK1AWYyD0jC5Ml/JAb3iIqzRfo8ORJsS3aGVBfHCL03Q5lz
cAe5AqVGOXc8NOlDHn745MRcupCRzJGSQreyQKHY1pbWyE4L7AupuXdxaanetykn
LgTOGN0mUBD35/CokbgBguq0h79jsHArYsIBWGz+IPM+9QsMkRm6iIsjFuwEMETB
8qg9WtOIs5iT35cz4mF8Sh9na1I1uKiAvIj4adDRkiXkLFp0Q03eZLQUEq3QHJyx
ea3yWaiyRT6OLnm+mCYPoDMNkSYJ3YxFQ2nU7ZmEvbIoC+wwgASsL7R/D/HlV/cG
syw17nxARJM3zxhAiKdAFN8TlMubxbTGvR76FVZTuyyJ1tO3Dq1K/l7gepq185yf
4sB1nGEChaHRlnLheEVp7xFkTXMn47joLuQYo8rdRwu7p/3PN17Jl7hKge9pYe7v
jFz1d+ut5ZUD3dotEeiZG3Q8U1ZXsyUsoY07v2QsZRgiJN6xaD/4yt6nxu2bBafF
l6+qm+GxlpvlzorE7k0Nx7IZYa1sDvf6sfupHg8MSZ3Yf+x1V8fgw5mZFYWSgGBJ
p6iavXB+wUwLKlXJ+yYXrlXjQ3EK8EhWhuOAVwQ0xBCTkLtxAc7D0ffaYMD4bwE/
2Ut4Dvvlf8V+gXOlo264orPA93NZGvByMbJ1fzv/6Yk4ntSEO9Hky1hf8ZtvbLNz
lTvco5CNWXaJHkp7Ji+3wniM6hX/ozoZcyYW7x9XCOWdiOXvx0oFQM3wT6GDL0ZH
Oz7VAbfyeexBwRiY8gAXbcz377ge51rEzrfE02uYY33PQ4JfLzOvKhXJwi27zp6G
/VuSxHustNUlEIQyHs5GoMvVIxqwG+7fO6IR1f2ffLkjW1PwiSrW+8Yzu7SWdFEr
TMPeB6h8IuCb8gLdIEgFRFaEBENChe3khQZhij98+u9F2UQBxFmuNiicUfDAfTx4
f1bZJ2FhXMNqPd0A5zGZfDd3EzNhIanrCFZbpE99KsAWN9F3QuPIpx840DvPkXJu
A0Bga2CAFiIgmgNoj34JiZ2LA7pKWTTTd+cM3OE+K3T7UJpESAfK7/YihL9rIqsA
51NRlSA8zauQz8tpqNpIQ4dNMNNg5bzQmxytK5AYed1US5s3esOPvxHEh3KKCLHu
B7M268ooMKehISvMVW900KolsCjg5AAtMHqDtvHBsYFXqUroxocyoyfTXyw1uAxr
aXgKBuFSXYNxBPPl5zEhLVweCN8vl++gCouIT0T1/cnmFUHCd6xddOX7qqFt6PhT
/O72qxaBZyN8f5MdavdSL/dPZwU3UEbcURJ20UyG2Md1JNgQFHbeOw5qSa3JsaPz
Gsgos6n6HQMxQN+ERTMfuDuNHGFhmJWkTO5ocbUKsVu/vksDMgml8WC7EiSFIjn9
uuSBgXJ9OMuGeOkiTXGxldtdppw7vD3rLjWJZJrXZlAXRdgEAAin61TTD0k7nJbp
IntnkLjfqdTFfOAmRpAMAgqH9KMxFqMNMDnq32a00gaInq8asq/0fXnmfPuBABeH
Ojbwk2KpbGzZHMmhedISEnK7CdCDRaVSBft03u/186HwbT8PR9hhPJoV9fexjkTs
mjGMR6WI0LtMqnDz6q43r+vlwuQyVOwfHcJqTaHe+c/aVfpk38eC/Yt/2jZ687vu
NsFjYDyo1mTV1/Bu/Mt6vNfQQYZgzjxXsv2P/lDnMNPcz9Aih48oy6GAkZ3Ipgel
5eR+uQbrmMP5HrhjhA20T9YVbm3jKs9sdiZ52Mzmvp5xnBY1XudKXv/Gp75UVm5N
8S/veWu6fLNTgg8zccVNPb9nZTglDj31cHHu82LFeHPK6B3377ze7YxX9FoHgGtu
2ON2JZom4AcKeFOYBB9IWzNcv2UTKNN8NqyaKMLnWQe4z8FS5tlz0vXJE0R0oNet
q4gONkEjFqdX2dzMqNg+F+6OfZ3TrOLSWSFzb8aPMhkT5lYGmYk8mpvwcThSRmqc
biNG9YFTceF2pv/Yhn3EihTEuJ5KUp1FikJWU7jF+T96zMibwaXwsD+Tq1YTQtk7
YB5qAkcSCwltYD8CIvTYfj89QhfA80EJq2DkRaE97/7pZ+HcOX4rLO846+slBCRE
GMGM8uzkibdax70PYLA7LbdOvhGMIa3hJGOLGen5hbQ+3Oaf88xFrNm6E48U+5Lg
/CB/24BjZ+orh+/WZChFbisJtfykMOEUsrIJE2LIJtixgRtZuRNXVfsBosmYOKbX
qZniw+rI+WoGGcRx3oofRjKipxoP0sLq7+/OCBCIjVVKih3P58NCbE2uWCZJz5X0
k0tuB6pQSuFBKjnpxSGJT4BKes6TcMLDzJYuejk+Z5SHiWHcdoikGhW23cTfM5wA
CqDE6ni8/aqmrGnc0unvvlfy/hdP0Pn+fsu64EnJd/DyE/4XjFiEpPWnBQ6fPs9f
O0dNMEVxsSd2RjE2AL7QyCsS4aoCc2EjQGiWeOcRFxih52KsGdIpvXAbH43asQAG
Q0LPyrKq+J5u6rXBQ26811PRvm5odO26pQHhW2y1nVQMH+0eBS1fb6B0F2KVCJ0I
e6E7dqscBcF/I6XF9qkLzBRyZS3H7bl7zV0lGQiQBsCb1ywXabqMilJvUfMzg/Ii
66EvNwnNizfBOROt+/CTmGg3rilfYzXb5AEFZGVJ8xGCvdZCxG+LIMTFQQjLasdb
Y0eoT+CvMMS7V/Kd90k8GXtxNV9VVITqQDYyOPbuaD7FNZMoZWO0Hgv+3NMYpcw/
4gIqu1yXvuytYY2Dm0ppkUHF9IJccLlKyslkVRVWd1QSLtfEg6U0TEKdMkQAgVp3
Lppf0FA6rypwpcAAlZVw7AiBOtT6387RDVi2vNCDvmFKgrFkBZU8ZHtPSqAOY6jr
ABlsIvEMcm5Ct816jV4GexTzRXd7mX6pJVkQwvqRLEm5h4shS92JfPwYaaq3N4tw
ixtId0HFWBDcnaXCN1j/GyFfctxshSasB4qcLPA0lu419dPDVDv8wRI8c8d/zolB
+b1nYronnc/afm48ele7oXmYE24z2Vr5fRTDE/o9+8XAUd793PI9XrpvpwgMslhT
rbQN+vjjQ7/Q0VTWhPD+6uLyulHYO1oWmsfNTqJRjBf1r0F9o7CEdkDiSeOqux+w
7wdXC8kW4tOTKXFH9VBYLA/O9hU7Oq6ZnXtH4EVLHNzooNsQ6mSgqLuemlo7Esko
vimse+N7aZN1jYzGGEZ0mxlM28wYW1u+QooLOJEfMG7Y3G89sDSMqfyb/K1jZZfY
ENJHi1dv3HfoBKflyaT2ZHUtTItb2m++TvZ7jBl12M00TdCyitTcxBZ74PbydU/e
3Xiv8XNoTEFbE9N11yaMJPb/2gY4U4ItEeg1s4bqRDwBBrxP7hF/S0s1CSqXj49i
lTyZmy/7rzKKWwfTJbrpOR1G+yiPIshhYtwUes90APHaIPpNUpzYf32M2FpCKMCY
TNnSCaQJNKPrV7M/xDNmQQIAQSiKCEHPP9kcYb4Bnnx0sSPJ5DJc84E3U3w2EGf5
SUYU1l1MHaBl4x/fcfevRw1J79Ou7y3ANk2ngnaqpsz/nWviZMIDlnAKvmkK40cW
Ai5103v5ZQ7f8G00IjxH3E1QsGK46gT0X8CjwesD2ZtxHQTNuk8BYz7I/d8sDtsk
BUEI+hMiJ8bd8c72b1k/Ql3EOFyB0vWrbtDJQzBtKLY7bCMFlbT9GwMJbXGlm8f6
YOPQT6fwAotXONvLtNJbG2yz8fHmm6F+X5N8t4T9YZ1tC8buChq8HusHcWFedRCl
E5+xeDjODqE6+IEVepmyI+mW0W52AZzJoJAztU9sXqpxu+Bi0dzuoOa1Yau9P7xJ
vghmVreODBeEeN19aAVhmJ6Zt/D0JrOSXiJLRjaK7reoZFA5EJJTdMUtmRSPtmTt
ilEGWZBJ3xH4Slu7pdJaNQjC4Vuz07hMW+ftKFknIYXQOwK+3fapmzOBxMo9eLyH
YReaIv0rk8Ami5z+mlACA4Csr534/U4INeLjvzf1rrqZXBL0gAVf2IOTjLQV/ehv
a9VyytREPpWF6tQWMNtaUi+9Rxvd04KbdbXugulvmOfcTk5G8LsULa2nSs76Vt6p
MyWepgcp+i2Qkj/evuKlE6iF0IGD1m4bcTL+3ZATRFaKtFueJBHdwGLJ/Sm/hL7l
TzTw6a8WbwwdFbPnBr5gKrozF7y01LeVZ5ErS5TPVXrHVgDEHZ9icCeJsPIL4QFG
WvKYlcWhBQK5GbGgduaUAvYB53MYUCOytBq/TKYHWDtcJnNDNxxtqKLLR0BxRg5d
T9DEDOkGhIfMi08kQ3DSKtIuTKrT3oHkNnaOh6en0TWsR2cqUg2ZNXjK9joGUmLV
0w+DD1gLPz5F9kcg6plb+qNkEkn44Mx8qjgfWYVm8bm7WEniboCsnobNvt+RCla/
WKmyoZciRvnVoXaXdVNbstO1gb7/479EMMzhzxcB/y854qF0IdJrjxL3bouLZU8y
hcXEj8EoM/kEAQL2hkE+q5js60daxZ6oCM4FHDvGsEIjepZfoOQ1I0W2GuIxAVxU
qHAv5t7hEuBdfi1r3FalTfHZHkVOSuzVSpbhcVC60DJPJH+lAVTGz7K5FFNNQC+6
2bd3f8/oiQUq4QnLMXjiwvroM7KZMYfZ6EcUF0dBedVxl6dAm9a+oGGOE9fVrf4u
w4jA4CmIMlUjcaNZ654GmLO9GggZmSqn132mlyze04aFCoXSu2dP5Jf1DVi0KZQE
aQmiKnyrsVyELt02eLrwLQNdAAw7aCA+0Me93gnaf8eIZjwfi/1YMvglGBSeTtWu
LuOfBks8K78v+VyCgT0oOrNU3n4lELz3ZDqsA4nXCApAiZKNJtfAeRo5bv092NRi
n+hHoqr4Kbo0wfPkEcbMLPsIKVobnf4ntBbjHuJo0oHDCk3BrwOavbspfXaid8aK
uzop0J2WuWIkAm7eq4RnmLTrteZ9H1ZUADkvOx9Q4y1otzBmebJtDyMbLsXS+lfL
Df0SCHdAC2XayzMiuIKb8VTesDbKtiBFnyO90GuHBKM2+twfCKWWZ1PGV3J9VBCz
y3p+WjsQjM/pDwte+HaPALzMUJ8hQkYjhD0pEeGfPdpHdyY/0OWCS1HqqnpGqisN
fJHP9FzzFpn/ZvHsKdUpI75s1liIuqSonaNlMU0AwJXgld+hlRCBfAJNa+qN9x+4
7zdDvktdBiY4ysEBwnli9UhNtcGt7Y11FzQxL38TxzE/b4whb8qlk/mGeNv4e+t7
43bgpQ03lefzO/7W4p9x7CP0s6dzD9Sn8FvacsqQQD7xCG5cICLyMRbEloHBNgBN
3T1axMuyQO/4Jc8ydzj/MvNOi0pl97L2IMQWbK69FitMXXsEfItc4g68IK42Okai
aGyBi6NxKyIkSpZNVRLXWrzYiqpCEfJA4I75pKZYT4cG/do/Faa1oKedDLb0uhFZ
cym8IJaxl/DTJz49Yf4aU4gmyraytXmF6gRUEmd+yOYIFpV21Uk3vq/LJJYv3PHy
dPMoCDR4SJoiJ8RHJfPJloBx0Z9ZTN63pmZmPuOzRVHTxF9RD5tvZSaLY+0U4kNv
lkGr6mrUjoF0nOZMnnWBkbSPGoh4ypHRWsMv8kFtbbsi3W1qu6moJDLwSAskFYqN
gJ2dApE+GP3F2spixMeoKxD6Ng3O5XO4v5cmhalk+HnAHmx4ON4lXqG7Lb6GaaPG
RwtfYQN1bwbJT5jySK7F+88J8dmQBC87J59zEFws2b8lsp86YRoV7AfX5VS6K0GP
cPgUv9ADRiSehl13PB7ky2qwYbsMTCrEUTPOMJA6r9exANC1XbnKOI9qmdaHFfe8
2dfKXdBPnsVZr0YgfvwGNoAIMD5l1JzaH/e74DOPTHwI/32deJDzpgYERv/PnMJO
OJPnoUXZ+gm10/UvmdzxLOHIZ2nFEyWBuzjoDJIVy3pfg5mwXwzjYh5aVwEZpIDN
UxI4aQaOedpJUQRNuhwfmtKViAebLcuDL+p6mCBBqmfoE/v0Mu2YBt5DKS9jLMvY
4+NYC4mHW/h/kOMUOjP12W0jDdMBVEQ8rNkKV8X81bSsk9h+QIyHHS272rKEH5P1
uHB/w0p+48Ywu1HXaD2AUEvRjvqXYRQXGONp3EOPG2nRahv5ojt6QP7m250nOoZp
wT8L1tKAa+4TtQoIe2ndxsn05s3d1u+z6+E2PU3A/fnJ35abuGU50IbbYIaTkMXV
I0fz4oRMWcqRdetP72VG13EfdeSsvvS9auQCYemlIJU8vtTgwJFwV1iUCb3T6i6U
Uh1QW3U/6oiykGBGzYW2q84cEH9DkKR9h+5qqiw4JopS3psGDoDvRe5agR4Xf6w5
y4ZZo6Ear9tlzQgWeSN09MiXZf0ZVZiheZ7w6sSvlxQE0zSXc7MLzgxLTrj0kN9n
Iak9W4PdnwsWQb+UgFpylvGhjTxaefbM6Y+wuEg7MlkBobrYC/7iGxzpbk3pKYH/
axuKu3yuk/UIUsJ/SKJqxwA9Po1k1HDWW3ub4X+crCw4AXurMkebfxcaiYw9aw79
eyJKX08UthFqmyCLWFVar7KVBEWnGCc3DCe0fHC+MHVh0okFyWuYlxOM3uObEsnu
O/BNPJGdyFry/ckQKxkC+6djbONlaRDzn5l2MIW/nUfktuKFIyF+nABn9oYlxcSu
yPIbcZcloDxHN/txEmGTFlPIObLCTOII4p56D7KOvkkbRWe8XRwWz1mlgOIb2zNw
XE0FvlV/YOqlkvsKgCJJeVgZthlNCAAj2ImWLsYxXt4R+TBcoZ0nFttfrErxnj2L
ZjeqUPnXN2KwmKs2V2b/ulpV5LkuvDUFvaEvxz3q4OlKm0Q0cFT+2UP1OVU8kT6v
aponewrzZ7GynB1Wk5Cug44yHdfB5klS2oyhFjWZulPKF7uNpO5Qgw80uREli6nD
RS3wJBfggm1cyuLD9aeVfEgFojiIsVgyLHV2p0nf2AMyGMgfJvGsl6BS4w35Z+md
W096pigZIFHZCPy1uF6v7tCR7c0VeliebE0TSIfEWZVCaziIOdjzymUzJkMP10Pk
wHujzIk7DXDIZVptoekx2ej72xV6L5aFTirlGyUCgx3Ws2cinMJ6NN2MNL1GkNvv
L3/whkvXtFvm0O5+DkZIJ//7Z8H5WwQNYcJaEbnoMAS/Ea3QhMmMm+1IeJlsGOqT
fVuF58T5LPDjAJsD882CUOi6sxT72AVeZxDv7jKThrkI4ZcI6GYn1zkyF6Z1gnCt
7b1tCNOsI1kqzq+J+5lSWcyKud5umZO4eoQn/hVPiiTf+ZArIvLNkuPjDATxmJsK
NKmoYR6yRFllJ92MaiA5ACaSf2m29RNVsttyC1EqOosKb78dDQCvA/WIjUgEpj6l
JMj7z8AML06SXYy77cvCpYY9alJX4EvPY4xlWUlajZWLxofbgpGub/8I+ifqVGrn
bt1voPMesUiv/HypHBuhVe9HmReUKicPVTq38x0vpXPjWYhOpG44m8OFuZXfJGce
HgELzq9Xtvgm6jb4KSoxypIppUcvYBA8biGQ0R9on6jzyxd/UZBy2Fp4F9oVYAJa
HqfOQ5bD/K72HOy+HrvERhAbXxDwpjlFUdEcDwLL3gYmMKuYgFewZCp62X5ORxe/
Jgpa9W+dKp/fuSAn/7oJKfCZ088DvAOebsmZrMXVpGlfsfogLscgijVQ+DQlf41o
IA8NhJwj/2iTtabiDNnLGxK+5OKDNICgOOu7Y2CCcoang8DGvlGfykA+xGfZS+91
6TwhbYXLpAG1SC+gB6VEqmaU8+v6ZYTyLFN7JteLsBipXOABzgJ8458nsO75Lb6Q
vYngCWpVRqGUa/bs3TX+xVTsfDlAU38wz1oSbBYj9TYLalBhnbHVBkgwMymztFAz
GkrWjJQx/c2ONYS/l7Pasd9PiRNfpW0nrappiONLcfOKqsZUrtR1kWHDElJYRlXO
Gyol5W8ctE84E7sTXEI3ENlvKdWCpZK6llFZvoOphNAcRTAXF+QA+YkF7JwUkMU7
v2/9V+kdg9HyAw8wHjoRdH43HITEPERUwvNeIBvY2kF3+oCSBYRC4WJ5CjOClwht
be1+qSpAsxfcppfV7Btv/0eAYKXImZScOLc3N2EXd4gf+EVdbE7aclXyfgP+q/kL
sg/PAYCx8nKyG1S/LhUTI49E/4D61tocxYYqmXToNV6aFxldV0YXdroO/XzO+7pi
p4EWhzxkKCQYjiFAawDpJxmc3jSDZIROc3jTbM96YcyoUBIbdzKlqif+cIkhL2Z9
1AL9xD9pOe4Bp2BmOy75QMLb2E9GBtxjnLjoJg7jm8Isw8dwlAAN+Dvil5MYk6wr
HSkm2P+kzDyLlGED2sgfZsqiNZGpB9G1NZifd3/QxsJJk+3VjQpSlU4FzqxZ5w1C
0gdT00ePR2XAy6FS45PBFphd/EUjXV3mJwSGFmS4RfHgkMSMP7bjv753+xgo3tKa
tzDGvXXTb0ylG0CrL1RkFJx58Ro+hzZSy3Mzebr3TvAP85w6+agMYOeH4cByaPFw
XKU1aBXmPBjEJwevCAMaTUonGFU4ynml9OFmPNg3WGMNz5CsTZJpQrCqKJj/hcMz
JEX0Szc3zWm+6KMNFyZ99DDojVcnwtLDvZvw83sEopwH13FiqPtSGkBoskQ6yeop
HFxslRtuC0KeG7zptn/VHukogP0YpVrEf+brA5cGtElLsqmvfNnXY9jofFnAAbCf
1J4L1GN9qbx8beWrwuIf+Xz5Y/tewL6+bwZY+XeR/fX0jRy0j4V6Ij7VvObwkTS8
NENE/utAn3rOarycb3C8JW/xEnXcU5QYXpk8q4cPXuJxMe+7U8Km6382tOWkVaxc
n5GglZTwHQUZ6yiNufvb6Ict40YLDyzPCbmUuW8Nu+Qf+yDgUh0VKhHaHJJ50OR5
VhExS8+cyp1sij13TfZD/vh7LfKkbtZxKcQVUbPsD1Iq+k0RAOtBBocjOfo8swLg
LiONk4dIMgnzIyyzvkFIDUenmcog4+6Cx4+gPOD8Xib1l9n2doym4BatlWbZQgwV
/k6QUh0eZ/6c5TjWb8VlK1nnMtUhN9lWdJfJ+7hjqv0OrTX6LMxJPn9mwygepyH5
IspZykV6k8yQcyHcXrXz6F7qJqxPmQ+9zkR+t+rgxHMXdAq+TJAeWHmEj5wb+pOt
8ZiZXalPNxmkM6GlnJb6Z7Rq6d0nh4NnC17pHx1toPmbYCUYNS+8kAoLB2X6h3T/
R9wpypVHavWD9rYP82kVNyrCr7MKXv7a50IReDUlNLY6YL9SuMgaQHenPVxQXVRQ
VS66Uei7XiV88JaJfj9Mc0LaN5iq4YSbGFAZ7krxxR1j8OX6HcNzQOUuVfOM/cZH
Sr6Q+S2iS7pZRuOuJIQH96rwDq/9QMztugwLcPWY3qG0tVPn2i9P7OKUzgK3f/1J
bhSR4UuNzCbQIoi9U/+qSmlXZHyeGIxzWohwRw5CkeGZmnt2L93DRO57Gpp2jjd6
7LhiyXzEB3Ei2XAUqOX9CBAoxqQ1j9uuzHTePrd6hGA49kc31EtLt4SC/Q6/Us9d
AvAxA5VkgdDsJGMYlKJ18LKRezcu9y+1fGeY6JzBbNwFRKtfW1aUJ68/0v85ZBvN
CkvAVVbTFRyA8jbq5gEG1n4m+6TcAcjXYfYTPvQBsVNckcUtagauggn3rECa21De
mDcT9T1DwDCB8NLfaLnC2JKF05WPoFOP8H+UAf5PcpfZfBOFK+8M6SndB8EF59m4
ZqjoEsBvItqiqwLNLFRwmhf0IP58Q4TsK6Y1AvZ87qPTC2F+5OJvS+5QcVgh24mf
BEe6NFaV30K7BRdd3AqZGkl7mG9eKDv+yqUuA7dhoFc9n9QE4S1zOGD8mkNXzzWL
5HnfdISMZ7+oRXwDUrbElseEHuCB8pMWG2Su7tQJeUfRa2Q1FuwV2Azop+tp/M5e
Poe9ZRdEgombmE4BIMlMZszpt9N6Iysh8PvZni2KZRePec/nV5oJYWY7dYkVbmfy
gfhXNgbj/tWXc8D1QAA66LZcgdAtB0gEiO6Sy5EdeRKCjpUvt7WGgRpwlXo6yxTn
qxeRRu9Vw7Jc3QRHHhQpuqjCJm3p0B68307/y7A8x4EKMBA3UFZ4Jt+bWdvgv6hs
cDfWvH2qlbABhyPRwVA29468+MADe5TtRWMmUBAW18EMZpDTz07a3vEWBHE8jhXL
aUxSIrpWH66fpYa/SzMGjsTqHRdzACa3aiOa0W5apQ/aGVvubzULgWvTgUBPaD/h
agyA+MdvF9zm06ioYpqMyacYA/IGiaHAJk1AR6h+U1vertnTaTVLpm+A5hoe8Wx5
MikWeagarjUBZZf5pF0LwrIEhnwTYf+TaCvQTywb6G658bZE9rJWp3uvaxKt4Cl6
KpwZuh3zWcX+eDRDrpk1NgX2siNeSyODZcBRISgf34+mTWlCWWhWRlgRvFDn7dys
wgjK0i7Ew4/6EaZpKzU4Qg8QGS2IYYcP1RCipk+w9/l/itEoROWnvDcgDbs5umXL
n1E92Zcet/FTzVLjVlsGaDM5/rODu2oHrNzVRC9uYR3iHyFrezPPchKymWnUznRk
DerSVC6h8nz9EQV58ZEViw5rMyojHHeTvUZBULUNmHEQ/WBeChMGjnSiDsMIn07y
hWW28f69TMRJPbX/la9ifOH7yKEVBF4z56+2BeziEuo2Mf9J+aEb/qenCB3dZNSN
ccBXKqX5fugdAJaFa1wfrHLgJAbsTpfguCIFjkEp2j+SFlVoYEHoK4Jm8blZv0y8
fA4pUySAV7/vxEZmnMB48We5XyefFbIlv9OTIzxzGhVNFDq8c2W91KeAW1vr7X0b
5k+X3YedbhRbuii7Ksn7LWp8+zlwcLIFXhWGueyKBRXo1o50+zWQbk9OztvoeoGm
fGfzcX2DUdbiasjJafYRCiMp4gI3YjF4v7ihuF30OcR4/yUbD5UQZUxb/l6pJcw+
IipGPU5UJ9APUZOynlcC0K5RDFz3mBVPLbJwYUVhamVbBYPH7zrEDv57rBl8sv2j
r3fgbx2No4DMDdbWUXR7j5K6xO2B/8hWn+m/BHpZ9VJgjSQZuZJcc/nwDT76adSn
Tlke4y5AU9cOFx2aPyRFijavjGCwQf9cl5a/5QiarJzWUsqpWgjteK9Nl3LNU79V
3O7u8ngCel/6t6Oc1Aq66/zk0kPKbTjWu4ke0IFInODSjceNRX9w5RJDuwmN54Ua
5N/UkffOfeqzHpVq//gx9Nko4wVGAafPgZ91S643NkXlZjmaMn+k01xOmz1ZgVpp
w5r8U714tPt1hVK+/+0Vfdu+Xg6CbTgzuAmXqbhBjVBsyN8Nr33kPF/voFegAbeh
txoTLxNNGDv93E+X77IrJCakvXJkG7lqnhfbeLC51xEIcsehbZk3akcCfG0MWAZA
pl6z6Xq5B1g5kXi11iUTuKimZU56TTkzidFkf0odIsiDs/XLEyxraE1qMSL3fI5O
DhYtOIti5GGW4Cq9Dr8tGn5hciGEABRNknAbDBvSl8dWTglEBDS+3I6KrAD2s8Xm
VpzWCm/xjw2dmV2cpknLKFYGLQJZuneorXRKuXwT4UkY1KYhYAannTD5OnsiLvTY
uHDBfAMUkOk+csMIf8M64YLDB0yVKfChEpg8qslLUnY9mrx/p76yZx5GYqG3FKUg
+tGOabsAYrvCPGBudvqVNcuZ6zMAVZApgA/G4JOBuhTu84NPdUhGIAxLg8ol3anl
ekAFh6JJZW8FHINStN9wYRHaXBQJK1j7/bn1hGDexdmST7zR+zt6Dg8q0MjoJUnP
NZjEwIDWuEYM8kTE+g7UovSu2crIY4mxpZ3Qri2sfT0sd+YhEV/pX3IG5PNpGWyN
joodmr4j5+sHcdADf+j2Oh+LA+hvj9BGB2ZXslI779vyExjA6cZ9yzL+YlFAuZ7y
xvTaMcj2zNIpxKYxllBc5Bj8Vh7i8rUecbrR6GVKEbuQ2y6C/c+GRMzE/zITLWbz
1FsCGuKqZYwHuAFnq1ZirzIxoizjgB1XrvlUQ1NciChTep3O2dVmoJf6mYnT3Wfu
azZ7F4rjZ6PfiCB0n+2CijDVfuZmGjHQkwdBD9cPwx9GnBk00lDOwU2Afbke2X/K
P81t/R3f/iAx5Cm+5ayknKFhtzC6VFXy5FNPTMSJ8xbAUlaHJlxb73v+wL6DT/n5
nGVj8H7QCCDImIDZ8KN/3jFHiizrWUev0UArDgNFbFZgj0BDXg2FmLX1S3NoDL0h
VGSTI6uaiK1pjvR3LKaNd4tUR7RZjsFc6PI7Py3XBNQVPJeKQ249e4cUE5pqfrv8
3fFgioLzYh4yUXKwqNlDdL0ZYYlTJQ0KJOo+gosNlnPjP7hb/sHGdmsG3QiOWheX
2BhTB0Qi2jsbb0suHoUqZg0+pB9yDBPBz7O7X55uV+7g2qIvd6tham6xf3N5cBfm
HqmUyES8o+WNFn9MvXxJCUSnPw4lcJWPPgpmp3B69Zr/eiC6NGWwaJyi3dFzW6iL
uVDKjOj/TK10GxG3fE30VNeIKWjzvv/n7cvyKjE4A2gBuaGMleCs9EjkgYJcy/zS
alSZApnFXvEnX5pkYlUW7ntbMDAvWCpxKqKe0M0xOOkjAIkhucXQZwY1Xu7Pi2DH
gm1nQthOkpQZiAK/YIwAHOVZkmPUByIX/dpzBPd8/6k90GwO79Fy0onhwa9p+dXL
HkQgxTCf0go/N7jEJkz7t25qf6ff+1YD0JRpJjKXRu4CoHq8kNCq7avDNR/+P/uR
br/knKTDKPbo8jbiusWRVwjPfmvEMUivwJhbjox66qRqHLXNdPGWpCpSV5ujgPZA
JUtytAcCt0tdQ9l9FTlGNPoNt8Xt1MiYkKoOWlCxmrUQdp8uKVFc001qA1R1fnpy
HrToCxt1dlVDD8dUbIKWHMf2LEwQWPrLHhHP0+5En60A+Ur/c0W8o6ihgySoPiNF
4+Li2pp+UYcyl24Z6JBKdUAW1nU22HGBJZ2DG2WVI88aAK2lLXJymNB9pDwB2utq
RLnaw6LWec05CqMJJPeNLxoddVUETPMYGJSWeOcgdirzkt4hCUe6agupNE+2yFXy
MT/H3HPOG0kYTbq88DjleG1K2qm+MBVBDUyKmxfh/6Rk3i3coPTaPeSc/CEJva+y
9ApYMp4z2r6TnJF8wHDp7ALd+KuSRk6wxgg6m2o0JPAvaAe0BWnh4ROBLMUClu/H
+e/R0JLd0jhtnlA/spMEfRg8opRD72dvmXRAqjftOQpOeebTLKy24mifRA4EK5or
1SpiPJfOnjtAFlewxZewpXqXtlTwV5+cPckvfaigdrIc4t4f+hTFiJY6TCxsS3M4
HhCU4gq656/ABBBqjaVgPsgV5ThJ472q0emQQY882CQljGdN5SBT5ppS3Ja+7fuF
pJUSjm26CdVIn0kepWSet1unUwl9bob8SaoO8kQTWjdR2dM+UU1MxZ91gLvVDF4Q
mn4j3b5hdYScxA6nXFnQ6FoPp3rS2QY4mCumeCJ5jDlU2brnE53pV+dWlOP0vxTA
mIPMCKSgU2YtOWqwhtVb5kCvGcKs9mtY3p4l40tAEDKC9yuIjBzlE7a2kBHBXKFU
pbLtV2NBKVop5JZAzxaRSbbm0H8T4CDj71GA+RfqH3ABnyMFu2ewQoBKMp+dUS5i
GjUlypTbz9ixBlekvYI3lq2F1FjmjXHFGqjle2Nt2HCpQyQExA0oGbrtiKfHjf4t
wJBCuoCE/4K3DzPZHNZLPPXybshwTAsdh5Hwb1Mb0qLD9qsodN2tQaO1NoQhdwpa
luO/wWhm7lUUByyZ86C+V9MXMj9vgP1bSgKkWvteEMpcI8DoOcty0L6Un8635A3o
LisfOk7dp8YuVxGB/pM+W03GjNZuUiPifYkykNhJ0J6Q5wI6Zy+dNPRFTF+GsEOZ
IGcLFiiLbX6Qf/Ek2xj4N3JFmLyKePVA3pWt6eEzLMf1bGI3wrYDUJHeKgO4HVgr
sWNnMkvI4PZ8o6JA4H+97ztnrfYRqxXwPe9zNa4DmP2d3nk6teTnXsDeOmbfJFiK
mw4+C51yQCe5yAEGLvKJOQACKAbwXCrWPKZocfh1KguBg/3JEn1aLOpxbRaxQWzs
BeFjYfpTE7l99e1WKwVg8/MdAJjJGI1YFS+u8iEBsNp/nHOOejCY5PCDBJQiq54d
hmlU2Fek2WPaFwEq6jS1VQG9siH5M0Gh0aT0O/ej1tDVRwJjSTI2ENfn4CkJHRLP
B0UytkMCWwl5PFp06qM3F0sFpp1PCABgebIaDXeT2g9YEtz4yBpNK06IRDKXZ35E
toaNvHpXfdH6fbzTV7jY2LGUF3zUi97Lic2mo9msMfXgB7K/o0p97d/piMZkoxGS
BKoAmK2u6DHgnGB9WR20XfiMkGpyuJyOFEg5MOLOuYAY7hCw0pMwPRVXeTtHv+Ol
i1zClvWPWa31ysigAXeUtXG2EhCIfFZBlkmWIINQ6GUG4L0z5tglkahXr3LU1oZj
jCqDJPjY8MXhvZiRs54V4fVQPxIWQDKreRZJJaC9IpiZMffrSFKtfNguzVOL0mH3
8ThC2AGffKvVy8aUI2iJFdoi0GgjVof8aQCkDLQAJPUYKp+5haia4Y1LGmifXkU9
HWncmtLtA9JGZz1uG3bH5zDydIOXtrho2NBfZbJNK6RWmG14MCxVY4XMrAMq1Xjo
i8VhVPPGBvtqbkbRom3bJpqrx/yi5s3A7xIbVtZjWsEowU5gTIYCx8Ryzo5dHT5t
c9U7ezCa/oFDIJpZdigXBZAB3/fvwhnEU1CAfDdACYNFwX+RZ12N4oencuPyZOLQ
8cxH5dDNtkt0MJ9d7hRPAtjyi70uqxRKVYcSZiRrU3GeFtH0W1a8L6POteP6B4Bu
01nREcVIjTblxNRP71RUIHQCAlCD44Su/4lK09X0QfCuy87IFPZcc8cEk6QpQGHG
mYYg7wXKVanWOjk1SglgE5GdYo3zxatwx2KLPP2Xo2Ur8zXg5DccvC19aUT1ZguW
VQkKBMnCCQRY2o7mRl/HwVTzskcMs2TSrvUlrvenuPvGoIjpGFybmXbWKoJDYGKq
pUsFQuNuDRkmtzz/Os9HOTEdhMY1n7Oz6HSQ5PBScFq9AtKbnkFzIB8etEO3UrBU
PZtzAIw4sZHzl+PHPRthLSVFk1Puidtd84zpnws20p6LLcSjXxx+1IO+7Hr+A3le
HgHWgkXHA6Zmws3MVG9wWstldopxaXUDyXPV6JxorhDjB1nN5Ov9g2tmpuQdqhSz
v7LWQUMqsfib7jOIY729K9jAn/XC+w0s2wRxtVb+kAfgK1Vtk6OvjqV15djNKzGJ
vvFNAn+wPUD1txL5bOqBZotxA3lnauJW/gzJqEgs57teCdrKS2r3TJJ5VllAjH8C
VkP45GDu+9PEAwwKXkBxgtRniYEHPEgGy9p01RguK4fW9SnHC+351VJwP0NBzLcx
j7ljHETgmQxSMo3LVIgQclZfctUiO7zAbaC0dAngR5s0edt8/lcIdZXtPmJibHli
dcGywsAODO5Aek007mFR0+SF5o/mPb9Jjdj867/fPNblvM7UjSZb0h0wNpUgK87B
478XtxjT1sebDHQ/kmmgLcUGQr+G7ztEIh6OQpA79AYQUrjEfyk6RmdUR92H4RBs
rWJsDehszY8Lt0HiDKS/Ufq2UNmb5F9rVEctOYy3EynLvrqsbT3sa1CmI8WstMJR
fdZa/f+iGwd40Dh1YoKPLbZvM1YGLA2h5QB8t+pLir27TBM9QNa5fRrCleZqVc1m
bj3WPntbmHvedkmAIShhd+Ss9vxPt78eI/y8bwGNFeYUspf4UBN33qjzvlSsGkoC
pOJeM2TLEjWAyO4+zU22ifIwYJv5aUJX232YiDiyrty7hktOXG6YLj4YBJO2gjOp
UgcIFZbIScFYoqBR/jH0dgTNSjnh0SUiSPOReRmO9QZEQ6EKbp7PxQbpWFFchP3j
PuyVjJkoCVha0hv4vu11bzclOkAHI5zVp9wzla3KMHhBjTFgvLkjjMmJOIedHPI3
GmRZRsv4JbsK4puyrK4+HA8b9r5ehwG+MH/IomUFc24v34g5y17jWKF8QOcwppOP
dPeA8RXR+J3G6/xaS2H/xHJhQQGi546bRXGzRyk/MMSr2L+JaO4acy6C3DVVGkzc
NLzdQX7b6JiwGqfxR2sv03fI/h7ly+YJVrx+5MxcpWzy/qyPP9k391PilgxxYvVo
P8jpnC0OpK8ub2I+VcWgLwiSCP+UcA5AtD9X4S0ou51L6f3P9ZVJap4CsUJ6haZu
2qihqwDOOX6c54X3vs7zMTXlcNqRe3AhmIafpQ2pz1xMfxr0yvl8+zgKzrdXJ4kl
5uf4OSALeKxX0uNbpgQj/qfp0eYJIyefcNIO6FKLODoB7PPIS274GDiG8xvYO5d4
iRHAFbfCFK594buJbQIwa/+T2gl1KjsCWlOxSnQYxn6teR4mXku79KoXVnaD5XLY
1g3ev191JwKXtBzI/angDy9njeiqSKWf7DV2yd0DZ6tiOhuYDl2tN6RkqpxCGNAU
ukF/bbYgmPHzc5BXJlQ75YdcgS27reBRNiJ7edEpT5Wa2HH8+s62zgHU9BwyW1XU
SYSSu0V11izOUUT0n/z9onGbjJx2/K7inaSL5M9eo1qLyka5C2hg+pCryjqa3mqf
FNm6E+sMw7mjxbgNobDg1LOQ59ydznmV5f7pTZYhtJBYsE1d+RMlqjg2RK/hRm0L
fSTA4McXRfESKSabUjaol/FaYpueg7j6WSWACR9yLrHE5hKscfA3KAcvT5u3/SWi
q2/S/m8Xr7o3IeR6fRrf7jsyeKHrr10RCm475/GMIYx6Ai7m+qODQcECmmaRJVw+
xt6uZ2+2141R+MLZBLHZRgTpWUjoqbtFVKAp5/X3wHu63pohJBQz+sLzeDWI5tWH
Mmi0npDZ+5ON5cNSQ5SmnGRtLbKevtmSvyAIyRpFBU4LdsVSEUHehXk7V9033oX+
bD8X7N67bgCigLEFn0vx8MkC3FODPwf2BcigcTzlKOFpIVJ57S72fEWDgvbWtnje
JpYTjfw0k6mFzwCH11q1ebGBkW9FZJinRXQa5P4gJpTu6dHFxJk6Vq8rdKp4qdBj
uh1QGbhz8wlVqqxme+j2JZPCF1x7o8VtWvMD1vDHJDQBzq3Xkg86nKr5npn3GOT0
Y0NHjLrLs4oJxtxCQzdMmbPflztD9TbYeOVZP613QMgwHOXXkKAErHQygstqFvLA
YU2aANH0XW2DrRGzwQ5KrTvMZDTOtMZIANiVl70CYGlA8qlGY3714zWsPoL7/Vzl
i1XhrxazPjMXYuH+IHNJt5PQiuP6tB+o6g/QDBxWDanJTNwNkdgvequrTgCTawZy
B/Qp6WPPb0oWPx28D5RQ9hlBOscLDSipmtmmQVyEoUucmdX2Xyyuz8XZ2OleguQ7
1tXYLBTDxDKnLn/QozqBzIfEgowNrT7aIV9qWxOhzHiKfc27dRheuAz9S45I4qe6
gVZWeIHOIDDGz52waz9EgEJ3nLtedIMKYI/sYjrc6AsLt5ypyfS20o08GfzAOYPX
/y+IVr01SYU40ToJrg1kPW7WaF7KoCPIeIYXyvJS0RELRvSgvsac0B9ExXs3g8MR
BOqui+kZPNiwxC0yHmz3V1LrpmntXa0P0a3IoGtTwpyOUOpEhlPicWLbOO19Bzxk
Y/Bu0++7uQkdVon4FLjLHHvszwbtxHo1Rd1+wJHEP42nHV27SDlzZZRBBkFcNF6Y
EhLi39nRTfis4LORcYzgaXX39b/aGGNidZ1mM6/JgRNuY483Zm2GT9yxDunJTG7u
Eb8s2CFnJCvvBtmPqjQ/1w6m9Wq4Eou6ywayTOAdi2/1jvACOGl5lpvPjb/yObnb
pkcpKmiayafWN0z3cmfrRNJRwTnya2Fbqrif1XAxmPhQ5BmnNTbs2OOEwQXnpWOz
6F+oODxclv/b1UsjXidkDgEembYP8KQzm7wD67kZ/80AeZYTFHRjgdVQxA6HGN8G
Lj+1ug/NJ+yEzH+ASPEbguAHTwj7GxVm9b4P3hK7B+sA4wyR3FXzxtdCyozBPzn2
kIhUj35OQqy2LOGG24bm07sujBHVQjCMQqWjX07HcpNjPasfqE50D+lqsXPPUwR4
yO5yiE5MXHRYQegNdCdWWKMmHf99g589Un2tT4TL6OuXEIe70tcXwAtAbyORkvi0
4zlOL83RinzjaIiHSMrB8CoomVC1yMY8ljs76V1Xigt8hLm9uiKFetp+UWrGHCzl
ymOpdXiKb24PewPEENeYWySU/mKgu3CahS8TRqtAUWySDX7AX6FUMr/FxDo5Y7HN
epukRYGrcia3ZwY9UKVU1ohQTGb7hE8J3OP4CGDL3dPNkJCHkxcVahFe8JuWJ8Jw
HKZYd+4XUIcD31UlcdcwPkfUEdu8EtfAs7EHL56V2Bqx+RtNk+2H9G83er0oTaC0
Qh39iEGb/Pq6gEY4LAcdEUKxI3+APIxtk4/NIRTc4057mKgrKADlOR7rRAL7/ETa
VZUb/rI9HuVzaA+O6+3OsDCuerA2DLpb056IotSvbhVwooKAC+ja3leioFSUG8/s
/5Fk2AZAl7sbQufxHJZ7LpscjQRWHqMyHmNqj2FklShgWaj/bTfzPSXEKcjVwKUy
95f5GzUBdsHGu4W59p2NlTRz30PRkfKxd+WD5H+CxuRszIt9RRvTuM3XUOD/LeM3
u9pacCu7Cwj6X0nRkzJoeF9NEt7GHEUbEun9uVP+OJmTXbfDOYHSPMSLgmIJe7mW
UK14CPSOyKKWtT8DYqRU5vRAoC2AYCtLMt1uZpeU5D9j2P5j1sAnvfr71H5YnF+i
4JEmW9AD72/FdiOPcYzITjuzr8uelceShDQYaRMNnGVtVUmsgH9KhlKdRAE4I4fs
fQAr/KtA2NmMQMnaZgIrOngld1GTDWF5EIfHfe4s6B2oCkDqMEBTWqauIMxpgaLh
xgrFOWdVh7uYC6R5a8jkFNaxbogVQRNLCuHvgOcxcicx7PjojvGaUY3ERjRhbfJA
xGrfLICydkid47cQCk0A2bY+4Tv2Z8cwCDXWjG1asA7lfknbogXIXCjWVQH2fGCf
vRI4mSs7B5T3Sd9gXUhnCENT8RNZPYtJvR24PiEaSxxYN/XSnmU1Thd4APdktRUX
NvvqP1LinCJOV8MqJiBWwk9RLypvpvwgAZm7jTcXKRhhO0A+gwVajIchz5n0tIS6
C0u9tt19NPwVbKdaWLxDVC3TGHtU7jKg1IfC7nXS1A9F9ZiXv6ZMOTO1p78/soh2
JeOLUNAT/RZX3qUUKVLaMKbCF6dC7u+c4+MPqxnEWkZ6kpnb2KHoceFEgixFLU3T
Z/RJLFJ4OArUKlu0ztfAIOZyqcfvJHhqmQG8Wh+sVIZohZdyQq1o/ThjOwhM1XhQ
5sAIwcbOUQ7yT/tVg10sp0VrpYguXk4rqMNhguNPF1Y/Gb/tYcMheKII+ha07/Wx
qUeS8EnnLqu3zGiLGGoDxaaJ4nOnlP9L5Z9U69HsnU1zAI3jw0A5bjOXQufb9l3z
fsF4VKRp8lqMTLOxNkVY2gbL4+QS/aT1Hwr7QwRsq9qe/JHlnBzFRgRRM3VAXnT9
y0O2Qxa7u4hLDzzWwq2ns0q4vqCl7dUaRtupRr1Xc2vZgRgxMEl3ld4KdvqBHhEk
vNVKcJgy6+qLL91aJss3vk9h4s2cFxRWvPSgBE0Q8EaXQyJ9MW0M6DK7GnZgNcSV
KznB7HT9P5htQiyDmWH3Hit16rO6qjRLTXDmFRAhohKX1yAVkAHCxCZWWeYOq/Cp
HrCIewMbj8tGFTjAVw8FC1ZXa1d8xsaMLt+tBvpyR7lEjkhMTF75sFyxJU4WU4/X
CoocYdeM/9uUxd1NYQvE9UGa+/Ktfz/w/8HHSoQMBybONuG5FzfITjHaUCJ3Dw9d
Jp1zoEomU8Vuig2/HH20Z9SvDyJgZB5paziTcQfPB9AxxGYSRyuSLTaPgF7NfcZU
8AuJYrIIkIVMDMRqJNNAEJIUWLNhtiKAaoYoba8fY9Tnku9icyaG3vpsWj1jI9Pc
PiBqRRgD4pxRQQP6+rxVz/ka+IdnA9EqBcB+1x2l/phrrmvIkVBJJXuQNU7tnLwi
GgxD2sjvo0KaJ+IBat+5/M/VN/FjE+NirXD7cyH0Wfn716qabpa+KwgP9C9MfRQ8
8bnuY6ZnC7Q5MzpDrtg5ERpxynt8Q/IQy+vrRZXgu6980XyYPFieyeNycsQ6mV4+
03CkLKFjb8CWhaxoyuT6gxPpSmVTQ+/k5hvEwIQk9cBeL9PgPoxd3RpcEoP3SZnY
OSxNCuXqxqPENd0WiO7OtYrg/PUPrvR8qpbVKrpQb2f+40s1DE4EC4H7xLZtpffU
GDaRlpbRE2nEJptllHeqAeGstnlHZCHGGuQpBeG7OFJO8sKqBzBxkQbEplVSI7kh
`pragma protect end_protected
