// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:25:51 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rkh+++yMZKeftBV+//m+f61EgPy1ojPlI4JCRQLQAMKyak4AVTLwQWPiYAofIwku
1p2vq7ICAu7BiEgbeeVj4cOslD05vz9SoLsQqc0y5GRft5VU/DDQcftEKCVFToh/
apCVv8FZIY9JySrCwnadw7iaMFeN145nWRhd14S31pw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3152)
lWaTErg0B8ByQj7U22H8qbUrS8EOhczacK1aIQLhUltScmoS6LlyyVm5R8rl4e+e
jH7Wl//hk8qjzjlPZrT4Xxhc89Arac935z+e9dgbUyDEuGaonF/8tgj1PdnqxQ62
VR2yljK32LooauEIwtk9Oeyg6y2Ww9ZRuxqarmJmkk0BMn2gjCnP11AqNEkmAXQY
aXA9lRvcYmneiV2e746BFzaDylCzkdnY0C/N6o/dJnbTxKbOY9eb8oeK0XBW6eFg
JegMoCeexguJJr3vMYuy8+PVmzAU0XdKhcvpWBcj2FVOHZTy83SaA9jaRpMDCz0u
j66IDr1IXqTNctMkOWs367T1CxQWBYMdhJ9Vhv1Mc1+LOByok5d4o0NxypCy2R9G
AkPVSamgwOnEc8KH+xCFOYG4XjhLRvhlcY5IayjwquU1yO6IVhRl/cOYvjOG1ygp
LG1TrhTAvzx0YAOX5QPJyYjuL6k1CrV/zcO+Tw1L2K4Zq2maSJnE/86p19NjeCZU
sYCLrM5eXuXd8yzmjUk8ODfvK63XRA+9qTu3IKegiMW2KdHeNiZnjZBuUA1iOyCW
/b/P8cKk94cOD7lcmnRHjGcF0U5iFZKQcRgvz1xyw03AcQJPrn+sI7VecT4dZ3g/
mc5PsSVsWYDBfXnZHk+FeRZUZzIPx9QETdnt6vJ3YSE+gJe+myk2eN+QzQyriDtv
1e6V928MNYYNz7XiVZM6/sf23ULOnLBgBWOpwmbKAsjtjHepvAcL9PEVGFCds4eP
Sj1dId9nCJSyMwdXzsLNHhLW3b9oC8kBkUJmGXLF0QbCLzMVmnxbit0ugiE11B5d
b2xya6ZLmdtrUZaKwTbFAEPmGcBLvkn0tkhC7kAVvNnAMnnxBrPe14KBeUc2h2gO
LQGvc5cLNhQKRKaI+xi55a3MQBVLZZ1A6jGVozJFn5KQbAhBhuKn8KiAXzw1ZYKm
irJC9yDoWbwS0+lMBDEcRougnvHn/P9dsHzOV8RJ+YfTjscg6RA253vaVnyvTP7O
yjGSEpGkfZeSXXvV4P7r/xurGZcgOaawDly7NAlRWc4mG3TUwvwVmd5uan75KF/R
E/CrWXWqWt9yAipfE4VDI/2LztfIxpHg+GSHcSR8CS1bnD37JOXkOxLT0jnCJUP2
gyIW6Ntnb6GjMnTzf9WZuxByRpaEHtKn1Gih6bpwPeZFdG6LxYHBg4KCAwKKpgN+
I4CLKdIjm23cxhxIBdl3qpJKw96TgEA6fD/loEMLF3jZ5rwCnme+Sus3VGEdgcc/
awCCLpzGvwHg3oSqkzWxbGLrhrJHIgmwgWMD0J8Zhri30ljwe4lt5Usqew/p6XO+
RbkQmJyV1No8qyK4j3DIav/Jt7CpSVT/0RMkpMaXaCwKK5SnusgBhG8sT/zkD18e
jARtvn8U6uFbz/lwXCQqnDeBEDgU41uJujXo7YOSgkohZJzcBooZKZC7ipeahjYS
A9G6tKlaJ2HJ/XUAWAOTc0Tm54ayJotQ5O5MrMt/Vma1j0xb9XYnuz1JZ7kEo3Sh
gWDVWg7n5KzSHH9o4ThjswyqYaksAKDhmGx5RCOKVijlIPZOdQSuxciupwXQMvP2
RBPSubTGPdUrFi0s5WTyrITXoPtWB9cx/k5DgrIJ8VgPKosv7FlxDia0rY2ZhfGc
Ko0Fj3bdDVEH2u4m98/RjeiwUyMfClrBw0BDvS37sf9+pm+GaOz9S5FfJaa340fP
uCzmkZXO4xuR7C69Fzqgk/Ci6phdgggStqTnBL9086YgC3d88Vyao/ZVE9bMoMFQ
cHDJP4y+1J+HtRecr07k+D8ZbMlvQImeClcOYe5cKd0WE3yUi78jpmFuHp5onUVd
x6Rjm0qVAP249+NC5A5QLP5jogJiVdH+zYyXklbTzmwIuzw3mxB16lxBYNUDKgrJ
zYsOz+T3H9NHJtwhmrcrgI3WvB/Imh9JpYaZz2p7JaWXr5k0u28+qvb86v7gWcAv
6b24GKkZDEK5B3VcU8JwXbldDVohKvsyil1V0ZCxFqqVAc87Qa8TC94biczT6lJm
bun255GfPt91p96qiHqGWsJW2KWr9qbtoCHykf/6DbyQSHJqI+YA7vt0tfRsl5D3
IkBdNfb600azpueAK9TS1jf2uqfe7OiH54HnjJSe1wj8io4qTQPDD75bQ7MbeInl
8j2NqlQV0TU5Fta+JHd6R7YlCVSY8+A2VR8Fedlv6KXf5ZNHHeuoX6silIgITYNe
0snWaLl851YxetAKkr7HGES6MLHGZQAVIVl9sQfggDdpN0H/P8dRjqYvVLkyZa6l
0C2GyPg5KpDMRUuYeTyPhN8U/K8hsXpd0QQgR0sCfMgUmhS//DIwoRj+6OAHth5I
/G0Xb9PvGHBGzanxbJJs6cNK8cUGnOa0pkIjBNourVfol0L5nb3ZBrw3tTQzyRJB
rrDV0S4mIAnC6lHjNxe70zy4sSzKs+b4alDXhlkQ4Rro7Iax4WTPAedLKfcFv2xP
u8VD9LRtS2OEi7HKzP0O1/NYdbZD6qMufKrQJslHubTFjuUfaCK3QvreBuQIMAOB
R8RFEs5hjF6hAG7LY6By1kN7dQPVo3344pQ5Y+X9SdnTpcf1FPRa8S/lJ3CAB26z
SrQsKY4wQ4jA0efK3yI5HmuvHfP4OMvqviDxZlvZBPp/tbUbWHplIXmdrxDLhAG2
jatsc+AsO0gI8+WmPT0YcdsGWnoR4+r7SzbY+bc6C9g3NTorn4Gx5yFyRZ4hZhyx
t4xl3KOsiNuGsMkMsuUUuSoMwH+uZbxIFVK/kxgjpHpW7nDqkCC3zEPAmrLsjB3E
/oA6vvh/kbug1zZLyFIBIjzQi+ThqRAkwvyvmN66p1bKZhMJ7E4oMdpbGSVy7Je7
9EPMcPxpHVgDCiVSY1g24hevYh34EtQwFfki6P4VVBX5BWQkZpUA4H92xOnw535j
3JTHec7GIK6RfImFGXo1wZMMGxruHcrrxu+SCaOAol64SRH8gWFQpELB4MYinse8
1OcevTI0sl4U5Ky3QDmmnpmBWx6WTkWeqCwV9O3sAXF/6htBfZVZJvyMpiSFmQst
AJ6Mo3P+OHXGnMsxWeBwa3WSm5haSPR31ZDiceIcwPlBqEbBqyoaoHeDPK21syjt
SoeClAGn6pgFTi3ZpL4Fh/ZvETMCb0djJBovzwE8JZanGt5N/7HvR0ZGGpLF6qQa
nYGc1YAgksePX/twWPDkYCsQ6Xj+Pfh37V2J7BL0XA/Jhou6PeoRsgXvSJaCBP2X
JW/2wHP0WlXt4jD5wnpMkjFb8JupprNgVFJM2sqRb3Ca3ASm7tR4QYCxkYjx8N54
/GI+tEgqPz19HorflBRBKtcTrzETh+rO8veSR03ZAXViQDVdJY1RCwL2qjSKTu+A
+ygE/uIx7psSrLucXA5YA+a7WPNTgWKXL7IvCU/IVV+NtBYM0JHs6c6bJezBHOGe
qoGmQGr6LZQVedosyS8cGnDgYyNBGJzfRH/7hv/PcF7ZxCZvxLBvv5BPSwvfTft9
jIERK7tuixfAPOW4KlPp0wEuHZtKkhGaMRqVAn/ZXF371GJqkL/VGM/MVtMPjiIJ
7h7xMwB6VPiRG8V2M7bspekKfKkieM2UbsJfgFwnPV9PEyRThTMvXsuzF1dkdKmB
4CagZN0U9+CoyIYU9K3KrcgQRoCR/ze+ErTmPE/3UD+82MbmkNSlLY806iI6Wy4u
p1582Qo99CUVnLz317KrN9tenZVvf4u6QP28EivucYDK4Nmq9bRqcmxfxMVeQCLk
SpUcy9nWbqy2PZiGmmftcdakKk50zMWlxMkkSfXfmpTULQikHSEssa1Dl1xPv+Z/
tTv5l3FDyZekmhRQQ4Jm2rLOlHDVe6g567dosJ+E47phsXyIKK26Qr11L4G0KQQy
TZhTh2+tAbVYWfJQiU0RNsa9qHJwuGj8QaItQOh7Iwd8FNIOD5qrK66PA2eArsYM
vhDKD/eK/B6szzyvh/Qv57QVivEC6rzdNOUwvPo6T8BiP8DfiQM4PX6lJGrpXC4+
QQdz2kFFv7GLNa3Cahd88lCFnU9pDabqmDh91l41HunzhyG2S5v9rv3wedGEKUfd
Af2WoDqqohqFSuUB/VfckO+Ja7e+umvdfdDERAcFnE+mytnpMARegXrenE7pAcSe
76pAyM9OlMk/UTY0yXGuj+iQy55XVBMzAOAgfJlX/Ss=
`pragma protect end_protected
