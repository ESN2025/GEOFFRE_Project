// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:25:51 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
shekQK/q/aOTcVsNDBbKCBVoWaq7lQXEFJuv1LdcvHbmCXEnnN8F6/HBDkPnnhuS
OZcWKExgrOlXth3LiiBWt+IGrpTRZsEqpeCX6g9HQck39ULxLRF4thjZjgUzayCJ
YFITrGGtv6jR0EEUh2rnlhwA+SpWafsThp5gMTUgiJ4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42544)
iiUavWbaXQm8QpQpqkiNvamWEJI0LdwF1ZT/zD25lSEtb889fo1p6odpk2/HqJBw
9j4NZqmxvyP04E4fJeIfO715I4WaYUmibmrBQf/bCKLaF61XgLXBL5qJNxa1lLBU
+qYz63LzQ9YPwe6MK7CKM0/RNEiOj66/eDVyRR9y9TLWNQJvhVv6n2hlv2scTol3
kq23EuYXSTUJdMGPEbjzwWKsOyBi9sTrd4gU0iqYmnU/GY5RuIegkXfmgGdtOHsP
0CDn6C5P1jBwV0MD9rB2m3eQCuZukIhrpiAJz37BAZQ0i58/jFYZj3DTWvw1K2na
8z2yUXB3OlELVwkwAKLze8tbKtPdAfn8133MpmWVWq/8DI0NGaAfWKUUtEfkl8xG
jpOAKwWT4UCUFQaauyfkhJ+SncAw+tUZPCk9J6/JYeL4NZzVPPAx05G1+IY4Wn0w
63/tNymhS/7T7oiepzixSHOAKIlw+KPvnejSEkVBhzfcWSISTLqKJ8d6SFy4BO3f
kxVdRAt5G6v5zw3uLL8lxNF1zRzuqGKmCAW1hYyv9M8W6DCXGQS4Z3XEjPFqwJUW
saVJpiungUt4OcJ6fR5p+T1/PkF8Z6lvp/xeVWUAUP/vwlsBcfGj7KRApehv6hNb
uazjiM6aSUkNnfG/cY7wOQqMJY5RscuUOqrBDVlMeIfygv0r88kxbu+uLKO62Gdq
ZxXuQnDGqlw5lE8xUxYZiaWcPWd6POKIX9PQ/+MylIVHpilWhLU35ReUS38XTHaj
tdGnkCk3ZoNbxhNbWSdknX7pRFobpkM0YvaWFQFQbgwZcB2cNkkIDVaI5yQG6L9F
HcR0f+2asH8aWq5ZYwhVwO6cTC18hXcBFtMdkyjJxCQIrUBtANOL2E78DS41nuBr
2dPZH+8rzfsohSrlkWrtlQ1gnBvJxXJ4oeThGgV8GMztIvD/9p85wzT4EC4kqcJW
xrfj2Pb5LWTIPMuCBTr71lof5yhrzB1ylHUqdqOE221xX6AaaB+b294Leb/6b1by
fAu4ue3AlcvNFGiV8jvC12OOeh8ij6PB6oCNSaaVSfSwspQmjQ/MW2/s50zcyaX/
iy8boFJP+R+MQKjsBRITSUkFeucGMgUEg7XusxLWWsiW1FzSjBrZjRFzMtrUqVn2
Xk9abRByAxAKJT4N34hpS3H3YVMWLikPAK76ZScgNKWidpbUGbDxCBym7SsT7FIy
S7idlXWGQlUAkws/6ZZQVmvxWivDwaosPlQoI1gfsYQRIwa7d4/k9GE2TefY66qP
RjnhwNeJfWyW/Qu8jgCC05AyUi+MHkh7SVq1EUxPVG5rYcn5g3EyH+1OAHVkBU3t
mEQeChR5hCXySWEibXgK+fFeC3tDLRlQ0qAK5rnUD3lh2FPTB52VCez/54VKbVw6
f8Mrrf1Rds7OHLbcGZY8k0FBLWdjSYs3BsDfqpS1zDKWaSnJkXcKXSCSsAicO5r5
Q2Jfi+aLEY8eVYZrOkXmUiCwOJODjTftVbcGtqb3Q70O9SB/DDte+BST+VTDClyZ
vPPdcOWo/TJZkEwu1tOafeZjNh1rI61JgmC6iavseYysxsddG+YyvgKI59UwMGvS
HSZkxVwJex71JyN8NTcxqFK2iFtBZ5nJ1/I0JdEXZ2fAyEWBveyUNpz3o8U/e9m+
eyvas6Q2Af6mMusxU7ek8ujSaC4r6z/wx4GUCQSjih9EaetsTusXLuDdFJ2txeP1
0dxnx7EJL67+CMA+5bJ0UPjqKvSD7E2T+7vENDybU0s8Eh8AhdC56HS/qbBLHTwC
O4pGkZBlbhMe65XSsFZ3mgzElxBq9K8Kyjqd2si+kvsMIZc+p8X9bbIbLPR3T/wQ
/HzcFmnDXWt7JUpjExJTftDnsI4/GcAorG586TdynxXgSK9wEtlPUBaUleudtTgd
AjuKSTe+G22USuv9Os+yebtwNZ5EXh7lA6ydvTgS4PY4L0FJ/tUEvGF0yABdnYg0
vIxbboggsKfq0M/ST7Pw5DI8vEkzuabrJQLtNl9TC7/tknPb6O6ao5r4R0vwfoIc
v8wKm4nqb8t+SHP4aR8ITjaP3A15C6B1lDBlAvL0jggsiSGzvT9hqKOCdM0dj3OK
lQu2d+f6RwdhYrXWeU8LvZpcHs8GlFJ/VUPljVIPuW3/2/ffDarD25MljSoKPmC7
c1Tkxls0y3JfxXzGEZVpIKBCIrEIwZ+5dgJaYAqRG1z4X8hDE52Yr3JyrorL7pP5
NqlKZvwKA6KsJiCM5sMzioT7JJ0Xh3C3VT9tm1b+hTFtG62ycvJmwEbKMRrlNUov
LzGALUQ1tIG7E/x6N3nu2DuFo/l14MDambur0gbO52u0GFl33LQFdFXtKeHr2lQs
UsvHxgm7tP9Dy4mxDxJy5jtzFkYTNsQ2PutTOYrCkmLg5MrQbVjis4lRcp7rZT+Z
fouFyMva4R1Q0lpiwl/SMpi8Vqc8CHKob0Tlsja5IXcLkx10Y8fy5CKmTus2gACM
3Keldkt6teZqf2uKZRxdJGLFCuyzIBgjVtqbtlGFyN2ErXTUS9MinejF4rXZQZpQ
ApaJ9/8F7tBbyNdAplXRSaoMDhvLuzt7K7Qx2Z56cHSWmKp9Ii6DgCykjitmJ7th
srD+hTVa3IAVvjtMYLmP9oYbjkUOFWqKAdN3eCqbH3z2XzElqu4L/8sccxTiSEz6
CPelSeP5Ui8FcwnA83y4jcjDi1+ety6VOYpv1ShZc9Ey4b50W8Tj4372GPvqZ0Jv
/A3RBFuNEKREj04ifrwOkKDkmy9hGCQipXHx9a0Ls0G1FXCg+U3A8nOba5Hc4og2
0/ihd64IHey69gdACc2U5P9OxKH3GNreneg0xF/wmmIoy6IAb7U0S014d3bb5co5
ZuvB59ZSFqoah0nygzlxphinNlz2zejmbCptCc2NxCrMWMF0Uwi7E+EM1l17PuBq
7vTccKK6pJZCI2lC4OS/exWzoPo3TS1u2MekMS4AHc3WG8bd9KdPdt6vQ8SkBSsH
Z93rHgtrqeoLThW/0YMW+lUTKnj6DicpPxNqCAtUHaM13RUWVfHvSyucgWHcFpgE
MoKa9y1cuBjggQMoCG6Bpwcf7Q156nfuamv0h4/ddJ9rK/Z+Fk6IUtZU540M0fqm
9X53q4+H7svYDju7IgtVJ2XJIrU5nFQW1cth9uv74vrfb7Yud3My5ts0RG79OxSl
6Ff1LB627HPpMCn4R5J8RwMzfWFZFtidjzIhzOSjwly3hsJrE89SmXKrBLd+/qdJ
y6YDLewsx+3OQ8Pdf7CQjBLxSCk0lJOLoqN6nkXEF6vQq5by+6JpbzjUAciMmo8k
YZkNqy/X0nErQ8y/WCEL0cpbDeqK6LwPLE3mv+++FJ/CZqx0bGmMmN4Nfnk16ynS
9qDnrP8z1+q4Entg9haZjYF/BVJqvyhCOz0zeDZLyilOXJ3/EVJMxNbYAUGySq/M
KfieOcn3zh0PBhy9MwDuDQPNDD6yK4yfViCGMKPQYta4Q7B02XI/Ut0ipL+psI+e
kPxSLEpWodvzFHOoVUKjKyIzgLneyS8pD8oS+fxf547lNwu7xQId8ztqf3yQv61V
EcVuxhrWg5KAQgYcN9+idm4II2QzAZFx9dxPOyw7s6jYdyF96EC43Da/SursUp90
0TnAi7InBcF5ITtPWaJIJRBetbT4ZZDdWmKR8QD1y0LnB5GUNJ/JvnpmfQGjNMcm
6fzHGGLvgnnIS3SW8/GEOW0/20pzZsdsUwArt6UcrWW7M1MBhzEAKDVH1y3cpI4F
WBLp/HvI0jkLfwSweLBPxhenH8SHQaEaKu6i9SAihgD5Pyd/ktSU4Bgk1reGtoXq
efghjhZLSBYDdVxzavqEHfRvBPjz8psezdWm6FW9YHDreKqSc6CNcVXtKnoxll/f
vCpscAmGc/BeLs8OG4OrFx7NGsRT9p8e4XdTLNSCfao2XBOM1LzVUUir9O699qPo
tVysUMD94g2hJ0VQCewxrJRr8nZcLhVtHaP0UykRNCIwRWxjz2e7wQzfc0yHh5m+
8ZXxfYujcJGRNPCUYrnw0HQSA8SV7PLvbfcV2j8mPi02f3cPgDXSbCao3qAXuEto
0FyhI1ExAo+lrEPk3ZwoVD122dfR4bAuGcNUI3wLwZ/CT6m7/n7aZS0LfGgNBG4d
c0ebvUkyBx3fhTuLQRBCz6E8N0T47PYDsT+LuW2Rah8Rk59PNpVa4tzb6CEkYEWl
a7TnYb+sATMVaPNTuFoJgFxWDnDeZ3wYPiMFSKYGd78xX+VSFbI1tWMloBNFrEc5
Rs+wFN+9Gl5DnsQTfV4v7sD4O5gFchAEAdPmEjvumopzGbnfjzoR7Jw2a2751UcL
p6UskV0xNnOWzCKSJEXx5dGMUSjylmpXXmx0sn/iuJKB22+RbTJOm2JIynI0grST
TJKUcgaYDI2TzX0v+YVXYH9Am8FAimPJ2mWq+dM6KRIZ1o6jNvCxbjdqW8grukED
2WGyk0Xqjr8JIxZOJ7c1iA01nXXQo3XBaiUQjqkCQC2pTMDpISut951QHIeUsHol
DpvsdnKkz1fjq7fiVjeB1UEjpGFZbh7G4CvIcuE/BWwv1lV3LWiJ9PFn3lp4leBj
7Gs6u/3F090cyUQntClM75aTJBO2MV/5MpMVBVgB5r8zt5zwwHuvJCpBuWO+F2VS
TNxkTtpa+qQDw9H/R1D78mGcqnnKaz2bFpZQohzqpaVt6HQaNxhyNeqO6K3uED4p
vQdy25nAtkoMejTSHHZ4jB+jbqxZhAm0JpASThyZ1HC2fQfB53RTs0Vob86drAgW
lg2oEkPHw3gkNOp5okRSMvBjLaRYS1BoE90MY5C5RcA5xnw/eqXCm1KTVSHtqGPG
RXWW0n3YfhVTRKqMJLR0n+ko4cLMIj+H9kX2H8nzRyQJ8+Rk5q5PEMSsC7TY/BMo
oSNK/wjNZaeOxHQNxw3blwuBl2uk35Yffp4K8gbwG/vdAQilZynnWWqskNf3Ofab
P++Rckddw+QcgfVZfSsqs+75hAvdDJYUgPHx7FoWNx0QNp5wlMtLFpbsqd42pJDI
PO4Jp4DSXao8cCWJQgNm42NW81O8t9iIS36rW0I5rrZb+J3+xunboTiMv3Vlr6rV
yYTj/6b6/gS9ns99rQ8qwPIQnpkgdpMUtkldmVcUQR5F2FoMIxvSZQ15vlwgSiVa
nkoUGYyuI2O2XV4h/txDABYGvkfhL7XzkTtJIEYR/Kx5/aLHf4p9VItSx0h7EueI
tGVU/d1zLSgEsp/HyxfC2TwVs1nwE0e/rgVScSqGvtU16LuS5gITIRq+OuSZ7qKX
X0EF2SHLwlzH2oJTFdXts3XFQAP7nZK9eynbLX9EINsmEzNMnBahH6JWnnraUqz8
BzH2iPIagoOoELrlcH+twIaDZKFJi/OMX4aqZlZz8tkdiMa98FseD+wY/0fq4bEQ
g/VgPkbd8PjYqB+iuWsjnm4XXf6WYVeob3jFciaYDdzTYUALJlkjymrdcXcIVQjJ
EsSNZpeXjc4eJoGQNjwP/vQI6GtyCz64pWr7o1DQLxnB4dSFoUaeg2Qz82xamfwf
Ufk1s4+Q5/NwmqC2II00gjRbhR36IHHLGj7j+E+a4weE0X0cJmsJ2LocHVmb1LlM
4+3NAI411k/pG7M4Awb0thbXbkghYzpAmJxfHLOQUvlgx0DHMcIKKnyXDCtu6JA3
q3KI2CJLiZDYSgq9SQPCFjQZ1iRIUKLPAyUW6vARCejSuEP78DD4pgtCndBBZKd+
EnQDhrvkCpIlq4ulCG3t17sQGMqxM94NyiZzXZdn7/ixW7bp3ikwKYD1bk4Ffy/n
da7fUGCbwPfbVfpD5BKOlJJDpLI7HOMPej99tglC4slsTCtPHmvjOvokFzrBzt8k
KhKFoZSVKMfe+RkuhqA68bUi2PR23YuCO9HuNk+saHaEFIWFCTo/x3J5TWqH3S67
N4B0Frg7ykB0mdsaO9/hUF1A2d7gnT5ZYJkbd+KkfVr2nEsgo6ePdP/kxWdQ+xn3
1SnAoaDKxAqWze0DvO7wLMuCKKeKq2cV/7+bZzZzuOKG6rcYzEGQHyBwC52aphkQ
jXN4/Ss07bgxVlauu9IDc2m6I7D0Gzt3kodrMGpL1GVFXR7BPMADZdjkBflWJXOm
Nl5qAMMzkzmLq0HurA55yfi6reomtFsAzhFJka/UwFCIm+M7CqndeY9I9MStECNp
AVY2uCT7X7Xc4WQM5uU/WIvohJCaMOKN7tkdXx2NOT32exWOx+m/OKs86rGwGaAP
M0k9fDyKDEFrF1efNhl46Ud9twtH7tAiTou2zu37C8JGRT5YL3Lsm5NVRkbdsIfE
8bbMubCX448W14CWzGp0nSWVJhxyRoveORadyI7sSW8C/xp9D3Sn1Z1R3/qLqQmM
6ttZqV+9R06zMLj5k4BCRCscQpIYzdxytciUP/1OzDqx5DQQf8x7H/tS++NCxyTE
FT9+9JTRgX0LaOqQnIiV1z3tLHVy44TZVIAGu7q4ZkntGSIz8VSmravTojbIIbc2
oKH27WNca1kZ4zgFwLVsnngajTJUcQQ8zYXgpQlAE86KagyIZwSg4XhGNXEkLLpf
rgJFUBDiqiUigITNHHwslrKR2aPMAyfLHBSMMsvIrRnsb/OIufk3XV0lLcPn3bIB
HfJtXnlAUMv1lym+59iVGxeM6d8qCOi1KN+MThGwGP1GGeiJx30lGE7X4Vxhfmpr
0z6S2JPjCrhf3H6wMgADeM9UAQMWFtXZ8iY5IxGPk9exsGuD7jSZGCU+TNtzFLp4
BPc9JAQHTgLj0TQo33xDxWPn1r4TtJUlxM1YskVUiIKdEFDLoBj2GtvDZg0i6RVN
1c0Y+TwnEL8fx3gk/s1nXKNqxmoYN8LUWuz/8Qo8kFvYNnrReS963WNTsHsFSTZO
6M+01pWt7F0dWKI0/Fd/zpm5yEFC0HT76vfK+bEazhNwSrgdiAvpho0cIlE8C2nS
+eZs5Ux+50iduzaTEZaNNFvgnlexipX35e0Fnfsi/YB7w5yLjLvgLej4rMAI7Isy
h0XkX/1Q53sR+0stjdMON7SbNESOCMv5UAx+n/PiLzdgir4MtvIE4PCo3xrWH19y
LKo1sH/NlUpmUr5oxPc4kw7qlu1rTq9WkuhNZlYAGSsa5JYj2D8FfWbkd4mDYXrA
/NUtBdb1Hxdd5dnH790Q4BaaxqeTWmKjnIv9xhpjdSIIeYNiIovd3O7l+yX/ulp7
bZpSg3gwOA706HTj6jHPDDjs8+a03ODHBZ0LqwuQ8mIh+pU86QhnJKHhmDC8UVyO
hDu9/aqsMxwlZjvXkO7nkFdOrZ6ABp8ZC67/tzgRQHRRXXDONq9fVWCoMlSDhgeg
mqB94OKALUbrxCAi3Zpwpgh61Vi1yOvLa1FK/wwk2hlBdXH9aFrikk77v3XtHq/U
opVm6CfTM2Scfau35OWsBraE5vNvf+K9NJa5uXO56qOVskjGaF48kHrBhIaf1yav
KYIJhOciElrP2bCakx4czddAORDT6BqstUutF8TEHqlTqTMept6otiG4ww86yeyX
hH16g5hlI0yWi44JVWB77O9/AC1JWh1JUJLwN3h3heMqTxUhPS7hnLqPoAG2wYCP
JTfCfartV0HSHa41CNTY/u/RjMTELxuE1RcEo/LTgtDnk0p9Jf6/e/H4x24Kvn3E
V2tjzcwzuPJQphhg2/uqv/cXoSkzqeZ8nlDPtTG3aiUwcaIth3+vto0vA6vKPlkZ
3cayxLt1e17V5vsgyZgT4NvLVS6t2Ej9T/ZVCO907BYjhYCMA0KAX1UlRZRBv8lK
gltplel4vlpMwF5lAeidecsVK2o+ybPSj7kLIzlifCVI/4GzADqpwaU6Vj+ei56P
jUxoFYuGh6ZxPlRTjYv8lw3iLRyTBSRz9RUVfx1r6SdO5TLTa2jmuIIXEyEvUdFK
AFHrSEa/1pN8KawN4X1kezm0i8anH61tCQLpwNAUcL5qCJcw3gxoJeKAADNwseET
+NitFxTMpmd5VZl/eJjf7R+vZe2Zuei7lu1866E5xKm7WFjIoRke32SLtdlTHpSp
VXrnNfHPrzjvDpmfRgPd5tKIXqjSnbVpbxZlIWuQWI0NL81hNOmS/jXtOxgqZM+y
QvYzvSAw6PpQhVOJGUXAhdTejwDpMNjvr9hJsuYlxP5d3aomCzbaik5AJEjX1Ad0
WUL8JejS38kuzyUvorknmy2bg7aAXF8hdKuwsYfZ5fcXo2fNhHrSM/jI1uYE/eCB
u9KEYny0QT1M2+611vakqMDG9B7ZdS6CiyIw0+N1/0FCnk66Soqwa+A+kP0o3CGA
A4voGMpULCJS8ODiSG5H+wkHD17ZacUYvBeG+IZ6WGg0jF5SsQMdgfQvTFbiHti6
3VlV+lqRkSC6kqIvxd/AKdWteXvahToOeG3fUYBC8gqjJOBihNivXztNrqYjlDV1
KC36dkrm8HFSHhE8OCDkXrBCNuYs8FDFVw3MHlTDl5NHU3cAF5lQ0YWWlltpgoXr
P+hX/P1wRkhBaWighTPL+5htHj8/lvnwx1XVgBvd2/D//oxxDyO2RXpJzhSH6LID
E24aG65zH6zASN17lN1auNCnkE7Nw7R+hOmGGZ/Y7PmLcF2tA/ds31TyoRvzDoK/
u7TyaTXMAIsUNM3zXYSNvo4dBXJjsYngb+Lb7vTcnPL554DBz8iCjuQhmV4IL6Cr
2Oh6oqAjGAVKvmHjFbfx7ABMirRGLAuwPqRHiJYmqdYgYYCk5oNUPciGgtpnhs+g
+3D962PUrSQX0JeaIuqxSInGJSg6yX3I+ZbzL0sp1/ID8njXtvoKgey8MwzLE635
NQDSeiR4kRU5SqduLA9obH1rRWdUHb0WAQn5dbwlHC8Bbk6rMDVoXj1iNvBpROUI
HW7e7S2EKYt9b5W4+2EZm7FUahzPny68Bi/2Cj8qnXCNttoYwNXoA9rMw3mhrzWc
hZJHditJLc4mkSUGnbM92eamK1iqE0cbl0s4CBXEj1IHRL09yCghTyL5WgTnEzsO
ihRh+/N7L9sQ8LmMqJrYh0RCCBgVt2EiuBxfOUcK33hhwRjwDIFmlHJB3JRJ7wri
XI+qh5CGxL4OmG2n0Th+JwZswB/3f1z6yokKtHa8pX1yRSoQ9Qar9lBrnEG/w7IB
EWYT9VItCTDov30Bfa/C7kqCEq7znSWA4r/F814Hp0TFQfDiuR+t5w9VtJCxU9m5
PwwQPU/DwYoWz5fH0c4dS82WtwSJJjLYx9PvGWgryaGeiIQ/j76+NSL+RO3bq9LB
hk5jYvL0xvuSU4xtmSwnZ/Q3feUbKfBJaRerwQ3NxKO9gyQeEj5QxMq9lNYcsVIm
wOBCLDU6IrQvatOK5+7/UCsFxudGHoxake1g8e/cVyqGvsJVZSpHO2afZhI1DbWP
LKm4QM8xBZp1RHIkmIpJwLr+XjEZor4fmnro9Y2fffytTJWPVFl3PTBtK7XMlRFd
yYKeVmIBR5TTsqfbXTckoAydTW7Q18+aeyWvb5kSMry8+GI/HQJHPOqroRl6IXT/
vmRSteU8C0QAj+WJjFouzI7lRfFTjdfYMkUyM+jpUqFRkjqf6c2HnoULVtdb3QGS
yv+b/RgKZCCkESTTCxI0grKBy1JuyaHhH7fQixZUu5zn3egX/clkCV2XOL5ZDlcE
beLbImyEMJx34l1GmNGzUF1lybal5chXME3lCJzw/uMfEU6yw6Ni+rWsIMGRh2GK
0UsTbKMkoqtVascRuiTHbxZo6We9FVI9os43lCcAEi7GzMCIhluIvZcqCI/BTLM0
/wNG97xcTUTa0UbbVZaCA8T1YYPSBhJfUNkH+9xNEjkIqF1pzQeTHXLppnRPi3DC
DzMYsWk9yTFS7XgOpGI9q2Ii3xvJYf4pfzjU4eGyPjkByJQZDjvvBaBGSLZOOHou
DE/6EgLcGBB9eDF2p2nwblMdRdvCxsGjvyZQk3z5ZVHyQbwEfyUNmayw0oXcAzPA
B7B2SV/ejmQ/aWrb3KpZIpAullVAws9+Lrt2Q90+uImEL9ekk5Hq2NKfobmtRvE7
bZaVApJ1xOZKo+n97vduUp8rZkRXJZrcbsZwWelh1XQXXNu4SzQdsR1i3nDIhdPn
lL19ViURVM7UssCgk9/1pt52+o2ov1XGoEjtXvO7wL3RGusE0C4xcJL1uotNc/E6
uLooBCG4AbZK6x2aeEE/hcjZHZU1zLa5tMZy4QP9QK1O/j2ZwtxDrv2BAMk2TMts
eC2aSVwL1mcYnbXHJx3g2jJW7vdMb2Ejgz7f1RDPHyw5WhBXV4o3XxdWGPVF3A+r
vj8LsewslJrUSY0csOm8Sm4GL/9QdaHkWmcRl9tqu5ABv03TBTkwBTNd+SJBGtMQ
99fY28MgpnbenW3JN4dtJs7ROrZBn96zJWxcLi74XihapOjd9YXBlGCqSiYHy0n2
WuFGdir1oz36Km+5akSXz9cRu7JHOMipEVxupM7DXdDC2PJVCXkpCUNpTDThdXta
sOqABEdiLZlBPpIo2b/Gvdxrn/YWyqPLiP18rx0OR3H9kFhEG3L+CZG6eQwcL69N
79izXbDIOwwRsD43CnuToqfE92sLo075gz/eRcU6FFWkb9QKZ8cPv7S/1TRsS0cn
W0aiwlbEoBd89kFZ5roni3MCP2MclK/4P+eEQMTnA7w2sIvAKQy/NT7mSh4ekPda
fZ97si+48VWnLxmvBoh8/k9IVv+Kcn06h/WK6kSsEbhC2Nx7WLkNtCM87cin2LfO
t8teLUxft7EQCK/jQRMTrVx/CZgfaJSD28hpQVa7jocKolAF9/pxIPDMLopuwJmE
tFBIOhNzfEwW4f68mSLQmoXDs1+mBS4sDwkKzTi18g8jsol+/AT9d9Bcf1dcB7Ux
27Cc/qywGmIiaF7y7ZnMbaZO8u4Q+BxyoE9B8zmQQzxjPrwVlkNF0C8B41J7ulkz
Tr3972BGzi+m9TMST2+jJmC64ZwC9tSq35hwBo/eJUYQ7j+upZvKhBSWqx2a4QfJ
FvDRTVAGso/dbQwuBZ1ZWii0aQnN7vTQ3dkkUBBtiztBHxFRIaRa8qYvfridgoyA
DHQecwcH/egpVVztHr1z3qJ4Q5z9hBR3xCw1m3Ujc+g/Jb0VfDSTy1lERPFYKWx2
DY+BOStO1S6xsxvzuFoQWHy4ZKvlnXAItsyWvMRSF6JcAWWUIGdelLkCOdymoZrX
5QhRpiKnpROiB3gqsB9noxZ2iPJQfSc1xLcFZGdFPuD8FqSPYB+1bLjRB9+oHxUN
xsCldLpiJDXKDdK8GRcQSV7fr+mOKyb6OuVo9x68zVRPXppCrgGF5tohN0n4/6Pu
dJtCoG8I1Or9dYzOXI1ViWTyLMmsqHbtR9SEc05Kkejr1JZg9RrfRrbMq9L2gTzY
PB1pcYad/mNkeFLcHg5NTZgaQ/+BrLBQniqw9yKZbfyRy05/gPK7urFPDuf6AIS1
JHF74+F5xDBku9YW6TgF/R2RNZiU/StBPChWHuUiZfK5pX3Wm6AXzhSMpMjGvcXf
ROmJ+dv1VkTi9gJmp2YIH6gogVa/oxID8+f7R0WdS2LfptbkS16gkgPs3WIw5Bls
SRasp+TY9pWw1iUMTJnc/zY6FueuoSbTnjnKkqOUeXDKvmRV9KlYRaHtTiTQYIpV
49a3l7/RjhZfzhbJ3rdl1SDasYv5IqVUOD7Vuhx2o2zUlt03X6ifNYA690t6Lgmp
qzRwuvSbhYNTAb0HAGzEqJryJi61CszRXwELaMwOMIZ9248B1Z1s0tI+5zTqxGPv
Rqzz0ZVTVpj2Eq6K67A+sAUWM5T+YPj5RRYN7eu7QlWc5j8Xpi0SK1ruVdeNcSEp
8YZWyP+NK3H5Rtue42yGnvkbkzoMDQa34tCjd5zs7PWPAygi1SveYDdALP+LmnXX
KmYQuMzQhpsig2ZuWBSfWbk3A+Uut8mOGWyRyBVNCDEIrCxStL7mk/G36WtCzAox
xdUCohy2ElpZYQmyr9gHg1BwMsvh8SAgtxX1ixQEBQJBZPMTu3mxeDUCDGjWdnUR
pgxjqZpBvg0/ybfcMvs3STU+6X5Q8YCYKmdTdW3mcMUWtfBUvM6/oWjFcXbuYo6y
12V+HrT7CSDUXvdtlbPdCtaZcTDjA2/Qa29/Rphm6PUeVeuaplWzVqA/uXdcFAfj
Ikkl/UbwRGKZml4f/dWGFU9SI6RJMjrtu7WCwZFFjKDZuyDO0ejAOTwvPGyC/slw
mCESTiI07gOhonEIKIrl4qKE9CzTctxtSPMp+Vr3L+SPdlMsfV9W883v3BOayVEr
tNemA+0na3fKTTSS1WCBZyoEVugdlJvjMrJASuGukuwkgsJsrttZIQsK8ynd3f3/
x9Nk2rDg10dzazQORBC6xkSuqYYxqo32P+FKZcUuA+Dw8uRidtQp+k4TkebO29Dd
cpIboiyygrdaqPuPHkGpKEpCRTKK5xuT5BExxqKBiGYZaMm2PkAHiW091rQFba8O
nSNGf4quOJfYWrwsT8tGNVOQhbKy2V/f4QNvDLc0MCXWkLdMVMMt5B+rJA141I0s
H+ZD1dtqGYszZhsotmxydfvtpNNttpTG6pQVSDRQ37syJrzcwflGfwy8YgdyoW1/
RAR0pbmWJqlEt5sjxd8t7rsB+fbJw/5yAct2SXFfLjkiuE/bnxrcl0g+qpBYgtkM
ZL3aGF7agp7vEK6alMW+NaZrK+fGOxsk7sN5O4K8uDt0jbptQI+dz1VeKOhtQ3tQ
zR1YFBHSO06YWWawI1DV9W/4qc3K1v2MqvMLTMIN0XxSeAZRggysWzThxJM9QwrA
V7cBKZ/0N+E8yzmoRgZEs6r42LQzgFr12DTGSH92xIJg3THe62OnskpjHnpbeEER
uiz7fpaZeKdv32Iuxfp1yN4RYpSXCGe6ty3pfsAsgHR3rsw0voF7yhEkbR/mj+It
uJQljqAgMfItxSiIO4DJaTo50Saqe7CrNzzVgtUrwZ876Ya8cmamVv21WzGN1oWV
eVsSsaU74I2UWAabXqYu9Y9Og5TJ5ry8URwb24owybzBbQ8bUs/sD7Ex+VKYvlKe
vYcYNELpMw4PO0uA96TwSn7F6HCPvFQWDGKVfo55pbM0zRUf7tvtg+zlVu+opLPm
EpqyAPnaVneZCstQbn+oqC8SxhSLhFozcF/d1QoaXGM55+iwhI7yDTOecFQpaDEf
1G2pSkU570+h9TJVswrTolIG/zIu9vbz4SwKC/14QAtZmrH9FggVBoxNEoAKi7hw
Q0kESm1BfBKl3ar0h0VGU6RlUofnwQWo5VDfI5Q05j1E6P7pPf0/Rr/TnPrCPLuH
dBcF1I/WGxS0cN9/8Ee1FKSNUjftoV8eXa1C2CRrf6Utek97nAb+NnjyE9EYUQDA
prDjTKn9kU5mjZcy4SvKYWhR+lRY2lNt529DnGLi26oblUT6TslzRjNt1J/QP5N0
2naCbEPR2wMmbygpIMkQnlNFQOBYw5o6bU+2G5y+qg0wEsc/boEaL5lT5ay8F3YL
8SguUgjmPwOouNcoH5sm7od0npEqWiw5B8Vp95NJ13ApIuwglL/AQOG9lmhOCh7T
bcTN6pi0wCvjdFB7MuooK7w8CiWfbRnzaqdZjIUKUvsU/srlM42fzXpqSwFZH4FT
Ce+Q0X6A0goBfKxDoBFrYgWM9HH7Oz4zMg9Gnc2zkNu1ECSgttF+WO9L2EpAQxc4
tnrm8n0S8Rq/ITeJa8RoxghLwbTPMgnf71e5WsIiSyw//VFdrJVFhRpALPaiqRG3
PbHFUQUarnv/mX3ohrwkj2RsQKiTh60jwFNW9ipoop6L18soCqBobIORK5CqPyIo
0tdarYj2ez4e2T+s8vrI9ka6hjldt2PONNS03N4AmYsreHwWPPJGoAPz6PLspIvu
hZ+gaKAH/2aDeDiLwNsLaa+dbjVH3dUYrm78PzxsNag5wdFRdscR7Mou2zlF47MZ
4/fCsxHreCtcbiS1OA/TuCTqU0Bx31p4QyfbivRXUltSKRQVL36nCWQB5A87856i
3Hq4dKGa5UmFoeIUmn5XFXpUhROfnK5x4cZUZE2+GeqO+ghzW1R9iFv5CV0Zd7q+
ZN0A5Fv6gNPfbSQ3xTntDEtrfvNPS683KS+ZYSNrG1Ph7EtNaHUYEcgWuVfRxtZL
OUFe8zIy8V6zATarNFVgR8djsgTpRfOxHahR0PN0n3XEt+BY9jSiPpPqC38AXO2T
nANvAOvT4a6yPsto3KOb6n5iDPhB0DwrLoXmVPSEqNhx1aPpYW0kD+3KqaNACUNM
TT4CCxtfelDx7/lylrjPyKsdkkpZa1IdhT5PycW5VT377fGE1fwgtbB++a1Dhykk
dqPIJI0uDX0Gpv8lbED+GwU3iopzarcnPqYVKBBswJ64SZ/B/BmNUb+csJnly5l3
0F0Uxe4LnCnN4HeKsiXCdshaMQzrFBFGCA0HxNrFycaq60xP3tAgdn2ZB1Y/rqs7
T2CRU5oeHYCLsAFWgdVoDlhItwMVXac2m+e2GojqSKlaE6m6zkBzncQsYqAO8ktB
QwzYkP3Q0FnHUN3nfbwvL5Kpe2VVYrgr5BRi6aOwbAmsysZIIEMgTQpMxvFlitzf
dfZXfs/YYkrxZW7IIXeLmMfCW1kFOxy5SDI3d2858I28aN+CCWM2bFPS3Nqwv25S
TF6y11gzI+887dolFcYliRrvdMTDmeiqnrt5GWcyUWvfNXDECPMsXcxhB6wgCn+P
tXETgfyoUgrJEZyZwe1j4iiz+yX13a4uG48ZArOMf50lc72XTBtUXazfctp/yoeC
493/6b+BJQ95wkdMU/8XNmG6oUmy7/+UWPHLSvbyLyIifZy2v4wDuVqDsWPwi53b
0QyPyZiXc5UMwD/4AXI7dzpEJQpQeHz6pZ6esylwH2lC6K+bITETS/daKGFzhM6s
byiIlNmJqL9xKbTqntBP1GjAlVvRWP2dcDXDfhmnXWIhWMlDhZ09LvbxEAwloYon
i9Lw3/YXcAHZFQa7dpp55eMuujBNzfzcUkUUbmjl4gOryk/5VvJ/zzIiQ/VbLq1h
RURV9hGjmlJlDlTWJdyHdmzHDf0pcoJ1vnUQvd0lLYtq2k/rH7uKat8nIdnTyPK7
Rv6N4Wi4uUPQrrOfhnTKO7wgwgUwl9t2sBygUpxB9AO01uQ8Xq0Ca6gwx3/b0+1p
PUrlu9BYkdvEs/+7BO023EMp7hzrRZ9bnjJ0t8Z5L2pc7zhFPrc9MjEqOT16b9DS
p9x+i5SmsFQjM3cEZC4TTailwGHcAsxuw6dLfSE0NaaLSfwt4sNaS7nRk727OjOC
IWOXLhhc1iGX1FuP4nDBce/AF+Cc8HHMicTzeV8XG62vz/QJBt6sSyRqQ6H0zYZu
r/+o5rxZHoX3O7/oJ9qD+0QDo0fCNKw4/b39Ds0DuleuYx5mpu/jcGTfWKPuQ74S
Ir5qVj5+sbGPuSIMJmmPLz0ANVeL8U/wrbtW2P8LeiMwYDoT4fYOlW1hMXu3y4wH
v6XjEITW/LCql6kaWSj/cQHZC+LFlfNv3gNEXyV9EG9gIoUKN8soDUzUkhhNpC3w
3/5G7IrZkXojhUQ2BgTfxPcW+LLNZDbftgYjx0z2+oJdTFr89zkqKjSb9bAtAJcZ
+hL27PMX0Qt5bbaF2XiynpV/WHk+VsrCErg08vSWdTiWV0DD6XG2oWK//m3qoFDq
+V7BXvDmJOCLSjffWAUkVx890xf15hIjTcmiPEglGiJWQT152m+U2WnMd0nCeDIr
tmzKlS9D2le/5lqM4bBBdhKMXZjlfZc3sMqa16YY1tuvxrcFd8L2q71mBNwlMEYr
NkTT2IrCEE1xDY5WzAnsySkF8KNBut6S2SDASubjYuuLUWbuDIAqdkKx3C/hWit1
zYmw2CBq0Hu+f9PNdktfG46cUVHztrlT18Mx5q3ImueWz71eAMX//zOF6Tr2qfFj
PUGh+BJG8xZwQOOR2e4KLNWCKSTi/GJZ8HjT4Nu7nHRP1AVoF24qA/qfbuOhD/4l
Jeyu0JgcYnnc0pZq3IO+Jztzw9RhGy2EAhJf+DUXlndp5FOsDOTork5gIPSuIobs
WGhm+cdWF2g7pO5AYcj7Ne00LLB91j7ISwikuMAzOG+zsht6bEbMgrs9tk2kQtL6
zhndmxNT6NGhVe28dRJP7qb5GGSiGOp7mVVjIzXcCyrJB1Ztp7faY/2ztY5LhGqP
a0bMzVoSQCVFSNicQjGYDcaTXc8NVf+pABoTPGQsVE+HcwSZHouIw4F/pHH8nZBR
e/m6H55uBjXitFjs+cd4FAFNdIjclbzTOe6j4TbI2pxQHtEHDPKWRFvHC+GUj6Pc
o67ytH49LA9tFuf6fQD39ySpfFx0OmqbJ67m0crDK8CMCrxmgSGttW0CnL3hh3Yo
cJSAeSl8drNtB/YMLn+lXPjTQ53VviVJJ6C03toe6WEo6nwn5Pi0puDkAQie/0O3
MsP8k1uxaMhE9VgsuCk3tY7+w6QdVNLxyoIT55OjNyAWghr3Pq9+V60Ov6b1q3ou
COkz6uEnMNfJVg23eYJBSdoF4TPnELzax/DOyZhMzrOXwnW2z1+FtqwloMxbTGDQ
E3tSulUgp6Sv+opqtM/8UVYKwIM11yi9vTueN3dSck8/ULB0NP/nJc/moZ/T9WgY
ymRaLH64eAua7/bLNRNHPyQWSdAAsakIwvwfny7p3LXGkknNf9P9sQ0+cAk77Hml
ZFu1dtVcFihikQn2di/o7nzgecDVNy+PPasnopI+LHcz4Ss/aTm0gs//8uwsKHoU
dAJu4HVNN5Xp25nV5jGwNJZkjcQlQ12KoGoCIRXZPgXfjJDhYZNwIitz3IUxzosC
N59wpvlPpBATrAu1q2yxckh014PanvigVaLn1pMFoDo8NZl7LULdfty5c2QjcHyk
Rf/GFFlPW+7hTPL1MN7+xgsOY+1Cfm2YZvKxvDbzZNPry7UKIREUbMZuLoORr6dc
ZwKTZjm4R6+8LzBBx/tOtJbWFv4B2fqxZCml9Eq5T4y1eaeqLAurvsNixpmSV9Zb
D6giXPQaxnOKwSkjn6At1jH2RZXVdnP0649rY8TQSRxRbWXIKs83mDFoX0+SWawr
WdL6mZxJCAEgBB66v4VKRhy5WtZpy1F+IzEDjV7d8CYklVS5JA1QIMuHLnAtekDv
iliFdjiPw1ClLn2D3Ym5dpflD7W5mvJ48uHkRTH1CbfXJdCkb+kqrBBZHOwqlUf3
gwdJD09pBEM2Exltb4hPLuybNdsH3vafVPHdPXIoKL6F/V8XjRMmYwxfyU0LaQiN
/KXLzblo6zl31Nhh8uhRNmIDjuboWZ/ADscb0AcxnlN03pZW+Xnzjy+Nrzgd6CCi
VucxylWInYjfwr5X+/KbIF35Wy/DIhuIkjP+AfwjQEEN91asR1b5V3HN9uzUKcXL
GcnTLUJ0TIXne+shGI+fiJ+GaxkvGtoDXXwNQbg003DhRB9k8s2cCIJ6pyrCjJS0
kTJA6Q0Pa387Ga0pRHWARhR0/ST9N+0ibbFL1cT+1JoZ2zgTS1RZ2vKHGBCABPd2
KAx76Q942LZXNxjsORI+n2J2V3boW5UtqRl+LZzCtsNBEX2tv6PfFQY23x60BFKQ
9DWBPXHbKx9pzRdey3vpSkgJU5ZsbFzu2jKsAGmxCkLiZcbjoLd20dB0H/BBA5q2
/CydcH9kZNKtQtPPZ2vEOSZm7rVoqwzMqm7aAMZL2vdqK3yHKrJaXb+zkmOLqaIn
A44TH7vwd2HL9kDW4gZVmN0QLpp1U9HHDYY2NBolna4m4HIvrRxr/tb/zg/7xrvx
7DsQ506MPAXnxG5HMs5mlbzYVUtcc5R5aB+WZwRWJMRP41UqeFmLW64gEqLFwGSz
WvfYWn9UyMrZiQBDAyAhd9ZG+qBNmKcxspwX53tf0h1fYwOCnW2RtDQY8hzhHfyD
6pIhHUcgsdHtOvNnSmaXZfQqd+wh1Waj2P/2oKDul/fYBq88jO3BGHHVyMHgnl2B
T4qirI6zH7aP75tR9upyg+uQmP95EcdxkHCcOR+XTYSC4/X/AYWhKyC3uZ1gL07p
nPG2l0ivoZyV8dr1HPS78RynswbfeDx9W7hPpmwzdV2hVs+W6LhsDOW1lImriHbi
vwyiiM+uwHqcD1P0UHSwJnrYBTdF6M+yF2Bzw7ML0fw/fvUbOueCNLBrfZdaQCib
8ShFRtM98XeJbz9QtS2CuvLWS8EftST/MWuR2oHiftHBaYViIg3RakKX4NKOSTSc
zkWyh/tppUugcZ8DBsaKqz10Nht1vcELX6WwjH3c8gqVVVq2PNijmvwERR74KRtk
A/EIvw6QOT8S9IV8uV/0qhXsI6N6r4wqQnKWoSTP/+Wqp4MJjdsGjuW+IDpEsA6t
FVFH3BwHjk+7zijozeJhFUarQUZ2SCdoTQ/8KZb0Nqew8NWcgEN0OK4oKRgW6qov
I51GfGkHn0vWXD1ctANwpwHTIVlWs/SydaZTrbaB8YLJjb3NYw7wiveMrCHGssq9
4ycauxwjpDcWNWT9tXsBvXzEU3tV8MsfCI0dkdDNHxr67wJaLYZ+MogbOT6K8sgA
Kb3oZ1NJOfkw+e3L0iHiIseaL+0iCgtF/b1kvyJsrY+X2wP2IPWKGeWVstofg45u
mYxn2/HZfuBkJssqxkf4zctHnQHisl4N211y8KkOB04QchTt81B7FcJ5mBy0+kZ7
EGVbL/qgHPOiDaELcwDIF4x3iOvnQQcqCIPrnncNWPG8NpaMLwNvrxe8/u7fXkwR
aMGo5RAMNQOyr4y+zrYhg1I9yy41m8WzMeOEqUZMcgrhmJZY79KIRJVSD4GsM0O1
T/Vjela9fNurPSAL/A0GhFzTi5DLdyuChMn9x3tJCXyQbUNzutNRfyCP02l4bCoW
ZFrrG7ZIQBqd1tfvs4DCtsrLr0iAipTP/SdWbi1Tr5zE/qLprUBrOu2aK871jOhL
stM14CijTpUAlCkcWaCaeUz2E2+NhnrXDEPuFRaPbvclDaAgSHzfAOnzvWxQnizQ
YCMaf2GpQvNx6W/mtZEOv7TSmjXZhObrr2losaP5JQQPJLrGwKv0T1BDYAC6AQyz
6Z8EHq/3Yr1wjSvRoW4GcntnMx+MOk+hJg93SprGg44OAh8g/aWX4Dn7INJ6jXj0
gJiamau5lrFlcFhCW1PorqDq9uUuautGe9Gl/hLhtF1qYmx6QFPz4WLA3oJaUgAs
M7YB+crllx+Lp0VoQCqPk8Uc06K31Ab9ES0ZkH3CapBJzU6gwypYQRTQfY3S5O7G
G8jFLwR8C1/VpEU6VN0xcbF22xH67kX6zUpK87MVaf/LPstYz3QyWcCoC4xUDajF
bMfH7v9Dp2oJLkAJw9oKqNDQQ46SauolFUiOIP5w9NBKAW1AAPsr7qp3izfL7sYT
Yt9Uxa5x76Lkra2r5wOGTWywy/I60rADpFy+/XdgKXxJUZ2a4K1X46g3XuQQ99Ud
W5xf51kHLG9MBxLk2p3DkKWqsMSgguzOY3vEsrarBwrJkGQjQcPA34+s9iCBb1VX
Mcf7qCCcqfJELmJ+tpzuDr+b4h/zCcQlskc0vLuMWVkxfbokLCbu1OgeQRMoy3HR
SAAZqzntSdGbwVwMknXz3vVFeaNCPNaYxVsCX8cStANKUl5C9vXdWf4q+fYAC1P2
X1RltsaSZ8TgCMUTSV/TR8Wuf3r/qweOMmp0NP+nmWIW+b18hDh5rSRhqL9m77wo
Z6xAxq8jrn2JUdhMez9grQFyooVypKFfeyv3FxsLVKYymy5cxyxUAcG/B41KNleJ
of4wu3BeQKNDwB5HJ0dBb63B9XqB3tIkdnNQPjrh8UrKqGsI6NDUxkXLM3HSpkd/
Ia9ECq5XWSh9fTiEG7B4El5+mJFhIK6Xf86eCsDw0S7EJmVWPZtmuimcUh2lQsl9
CLF0yp26H4nvAFMjM6DWJ78e9jNoRpHWe3czG5j5+qIecubhPSYb1xOzDPG3Wd78
rsL0cfPExfPIqDFFGffapiRFm0ftPc5R89THo6mmemHLX85UglDewVOCtsxucmNF
Qchn/nu2p1Uje2UKmbPi5U16E7KNlJi6Y+Otwl1VF24Zo5AId83R9walTDOCEFle
knaDE/VYm/v1nQROzSzblV2wwLnrP5jrL7wDqjK/jb5CYcAMTYXdAUmz4D8bZWnK
E9NcThegH00HnKvfI6TLrkx42iDLNsiyTJ30xRlyawC7P9uNtEBYT6ePHSFN+dRy
zHDwhQVTpkKoaW87tD5eNX/frhMQjh6T2DYdNEPRQWwzKsQgWK9aR+dIsckn0IuY
OF6Vg4oXEVWvUpfmyGtPjSsDxat3Fxk05/uEwh2+XmWf1IFzkE1w8josk/0LM2mD
ZU7Yp+DsPWDTt/hv/oqAvmwj9sCPIo0QBhZbBtzMA4uptt13iK+hNBJUXLWyULVD
ApQycJ35j/iAELM97Bp5qLWSpkPg+3u2z5mRHoqtMajUhzZNUlrOuJ9wDSAZB0+L
nLHsD4+OdQCrXBMeuMePZHograP6gDfaBBYbEdjOetutvxu62deOMcs/hcq2jTnk
lHNnPNilBD5lTJTL81GycB8C0mzSr2T22WyDUxgwYEH+hSw2uBFjFOw0IOfaRbXv
JDz5NFO/HTmsW5dX7oT8CgseY2EakQRBl0+EDaT8WS8yGDznqV7/Q1YUro8dXVOb
wC48LuDMih7e/nwovswd7UNk8p52uDi9w0dsD3T1NiO7jJ8UwHtsPl//a7du2RY8
7q38mNDjMZKmssnddH9z533gy1EAuh/vl2NNDLzBUEdIHFFizBn3JpopCiejguxC
gJy1kMn7Kd2N7aUDDire8LKUMcJ1Ja2muEdg6FeiVhkmao702+s8CL4J9L5UkOqM
H+47Sq5WLcihjO2yl7yQptix1zOVRxZQTJIukYqJV7rzatlCN95YdTSF3EUWGkZ4
V61Yf0dpRG3yjXfL7H7ZW/outXYOJXLwV2O5+gy2ETezE9Un9srF+k0FzG0Ot9e+
IanIDMDW865i6pBTpyX2/6XYO71NSJP2IlX4qTbMfgHVsXfTxERQLAHxNtxRCS6X
Aiv/htdM2VgfGtwPCY6N7zG0SRnj2N56xrunPKqp3YUNm7I4c32VOLtFIxXcHSrW
SBLtk9/2IQK62DH0HSmr1DX8kPrewjxN47jXn5ymZZCMj2FWxmoH2nr2OqgI1HJh
3e/k0z0thsdZsmnAqXZw+b0u3TLEo+R831Puhv2ENsPqqR+yQsjuzsIdH2pl9T2G
ghxAEFy9uhE/CHRSxWsk3MYKD1fL3hJ39KPV9s98eAN7wDpEcYSwdjyNLNdYeQD+
/iNxnUSz5gf2Fd3g9qyzvtJHV8fYZLsegHv4dp8I/W9ExiQvlUvu4FT2srsTw4GI
AmRlvpmXdzEQ1r8wUA6W8J1Iy0x8iBe6ACuvnAjCAJ8Q8rurkDDMnEP1Qt9S8XUU
8XD5T1K41Kf682JuxlGDP2sKfG7xQirFiIAcNjXhtqqHOV1Oj7p7M0+tWbw1h2iZ
hTeBJuWoPq3f3p/g/KN4q0v6Y8+bJQJddBnryyxP4R106JXfR5br435AXjrWJk9+
irgKHlB8/6objYOPCpCJ2fXVF5edMErG7jL3+8STPYjo9is5ehUtT3DKMzlEUu0d
8QtkKqG/bf7nyysBuoOiBUfYy5XGkLDcbtWKX85UykQ0orpVzB2hhUBKr/CJKBXB
nFslkoti1oT42Sozjgs6HhGcWgT1ADbDAjFVT8TGJF9LKujwtMQX8liWjh6hoY+f
0F2ulnRrT3v7rkmHyqkP+QFcBWbMEl6iCqshoxBjNRO1zef1k18Lnbxudpuw2mKI
+02G0rZtASWobTVmhcyvogJnav/77pwE+7BxbF26LHRE6r11T4tsSMJz/d7tw7Rb
f91HAk0zgpT7/xFKnAuk1dJh1cqeaZ3sJU65I79p8wG3Jno5jthMCC+mdbbKm5i7
f2ltzeXMQNr2uOsNweVYmCzlcdA+VSL/tKbLSC9/wnQ74woxcyqlcsWKyVIOzvBt
a2V4Fwe6iFtEFtUOowPXDUN6vhmQeX+FNziHNLRJBwMxdQLL7ocnkG6XdqFjblya
M+xjG6yWY6+DYZ5yELChO3Q1k/fgm4VuULZHS2ktVQyTAUFLh/1LNxbI0JliEPsL
NXFptJfZ7vqxqiyVnah0x8J67M1ltMJbGerFP6tkBa02gj7ComLxYiBECuzYL0Uk
EjAZYZBneS2xMmc2TpeOydPXCKx0cABE2kW7q0TCtvmlFwIGIZx1KWtzLlF/9aUa
qRmtgO8tBR7wV9TchLbTltFoveNqS+ORLUbP6DAyMO9RB/GF2Nu8eTBcexkpq4hz
RLtwvDZt2V/zN4WRd6OvVZ+SD7siiJoBoL5u2DQUJJgzagtr+vIj2P99MJKkvJIA
BvE3K5Uzi6MDZCXRYnNRrEstvDrIakHb2hAM27suW72CzneRkq//lzDpp7iovwId
1zcyx1742FTVKlaDh8J+HaD8VhyotgoqGbEVYg0p2hM2cn12KEompaaV9MuOMQoE
zZF4h0MtID057ZMGbomjMJZYmmXxL7hWjDWXWHhoTy2n6aHfsh+9eVD/i9k/SPWE
bASgUOD8H1/o/RiLKQ2rU7GlLb20yWMN9+MP2VkL/knioGZJNZE50p7P3HnlrKkZ
MwjD8Skf8dpBSZG7vf23CdYAi1yLbth5Sk5UfetX1elcn9zUTJh8e38xmcOA85x1
wtUcffayyBt1ur07wU8WV4GGbpwnWkbtJRtDip68nm3euE1P6h9nVdzWZhHUjssH
aPQKQpCVN9+9p/1vTG8PD4qwzuOkgWYM8qEQ1zVOX09J6+P3Fz8Iix7qx59uqNnr
gdp9LiFj+XQOY4TfSmXsxTYk5eaEwVv0hliGpfR6Kpy4LiGcTQcRXHVhHpkc6UlA
+77UDX1UXsaEImqD8BnWnyJcNGXqr5ygR6OXKl49Uho93pybVN+bCrtZ5KpmTnop
C5OQMueaudTTLtlT0UXw8zTVoHnwa19Nsj0wseh71W2RmqwVEjWdW0H1WvvA8fgV
wYquiNtVjJOLxtHwQwwwvLI4H00eVfU9iATuAXTcWYtfcR8bE1UtHm9NZCUnQ7nK
RehuYNWsd7bgh89AQ057U7C0TzCq8AGuftlQWs0Yjzs4PoiQMkiPEieIxP4JeYHC
H1EN/xaaOuMFvgJABygvE8h5vfR9qrjUoj/l2wFcEVv1lNYasyOYodgExHanI7hD
if78Dmz9JeicI9+I8Wp/OfLFCSSAiXgAKlZ3xG5V0HL41DpJOsOeaGJizwik62sX
d6pwMcG6eirQHWENbneFWwXDnFV3qTXkaySmKPtgmZOdhrW87Qy8sYvfsncR+KdG
+36nDNkQ4idNw5VMt7+QzzSqItodorS0xbjZEt+IHnZB91PpOcFKYNlOWxuOFxzK
eBWxL3Pe6Lc7jdcdEHFKoFvhmyUIFPbMLOKLhRgKaetwtjdYO81Bs0ia73zd26vg
3I/dYr9+4fcuub3liOruL6hGcp+uMbdv5u7GKt27nFG9vhz+h+18U6HTFPz1TeQA
sLhoya8n+MtLSp6CehCbmuTp1Cp605+IybJDpmBZP9XzBSR2FYUNOhaPI65gozYK
fFpoZLFkDBw5sdQ2ZyQgle/KPPgDf/VZzbZ8Tndnsrc+9gdoqNA8wqucztvD0WLW
v30QX9vRyJ7TNQHSyDnIkHqsen3oKs3Uc8zmiEXfbXsSGLo6bsJIN+FyytEFeLf5
ixWzsg2Wt0jRTwKJWvacaj99KeHcbzRRdd8DhzJ3PGZAj0gZkGOyRZVjSWEn8ke6
99zJ1/L/oeUhf6wUpGs0Q/t1AUSjefLhAPP9YGC931BoKilmtMAPGd1bGmBxypkH
uqLkogr+mjgmM2EEzUsT4pG6nDBVY1OA70ZTDbxSShAZuiNNjSHTZ6R/Q73yOc0O
p+fl9Z3c9XgH7o/8O+8mItmyRvff1AYQnxxCFnJ0QPyWLVMiu9yZeVNjuR9/R1E5
9HwQcFsCzDaB21XgRtxWXtp95QbaZMnSnxR9kN/ujbIhEvHSO0/ADvrJkVrTrB9x
nYqs6FdgPJAeOxhmmKDbQaAYWMVHIFajgwF5BUhvBdFkgrcfG4traXgOfPy7lb98
A0f+PjU8F4Ef4DsUCV0kkV4HGjQUEHH5n0kdH46OmHhLS6Id7NKJJohF3k4o5JO0
g+z4JOtOeqeJ6K53T8gcFjPPWbcM1aZkrJXwJTXnQIM9JDRqXfisc0W/zE33J+yu
CdR7sW9NEbetnnlfEmBSziz7BmGxVOLouCu52/SktsKkkp5PnDZSCnrKlL09NJDt
Os5nbmnAqoFdG6tB0R2yDqkFH+YOcaCe5sgRicyNNMOCo6qU1p8hlOwE954KaqmN
gicT3H6CQ+g9GeDSYkQ0cNNpcXPzvdqrmrdOkDZksR/bgPpvrMnnbdGfDjTN2sq/
1GrZpbV6WnugbWz98m6dHl48KwtIv9fs1/FYJjOrie73T1nkD4O98jrpsVe23ztP
iStBudf1z3NqJ1jlFkQz/iDwJuikIpT+5wkJZfKn2ciR7rKCodHmHmzAJpxk4Dy+
A6hGfv9fTkBZIwck/qh2aKHem66rZLzHzwWFy0ePmH8YBe0jTvDwT7tDI0wCEWqk
080oORnvNxU7oZtv12z6mIAbyxpctQGKZJDlA+hY4LzeaRFV59+ENfUreWmMeKfH
rK+1VG0Tm8Pmo+qgS1jXW6i40SOhZppAwI5hgQ015HrA9xsV8/K5CuOqPkm7yM3P
2OdlRxxInGqY5lt6v1oNOMhaHYbfF7Q7uouAT5L7ipOaV2lJSGCj0U1e69bMGLT6
uV1C1OhLDQFYQ7VegLasAL83j7aR7TS7AaOOIVvccA1Qq4aaDo0z4PNP2TL5tzeL
8marT0D51q3Wrn5I2QYe+Xz9uBwxmV59DieFSzKVN3d0+JR+V+fY5VHSX86aiAjO
5+KCU2r5+GUiGrao+p/J75FIg6+vgxKxRiZE7gZuCcEtQkDkdD4lto0GmczUJxnA
e3ra/FT29jBnHOrKzaRbplJtunxiOv8mIY+OjixddChZNnCHYWV5IJewxS/vtSVo
I40VUYleqoGhJ4FnvqZok935iuYtuFmy8aTcxZYmolIP4DCHbN0iONQDn6/86OY1
JrH4TLaGmI9rRAdpHVJVlVHUIhukY0VL4wfB7mQaDEg8c9iB0LXz6aKYLP5s1xLD
w5qyLAdCLjBSRuUSX/yMzXfhylhu05y4Xw8AIyMSwIR4G3psJXrEfwFowAWcAloG
+QyEqUn6KBaGkoT+w0vyvd9eaBOHoPNLVIyyxxCQByvfOCG84gZ01iWI8ROaZ2sp
BsWoIcKbc5d6aB4uPIS8KbS3iJupppYLkTG5mFSD0SnKPBlJo+g9oHRfN75reF/4
IsENnp6wr443rdRR3QdZj7i6W3N4n183GaY6rV4mwKfP0x+10p/GIM+tv4WdrnUs
Zbf82tBpywTHV8aF98Z3lcu4l80vjar5qKg/nfFTkQ9RemJtV0cYpCmiXE1LD7E5
m733LEy6KtugwoJPWCmr07fe8iLyrvpVlEY1QSB+xqVmoAs0X5gQz0i1udSu+mb0
FHnnDy9L87qN5QTbhypbSdCa/3bcuWhyy0iA8MlxBmouIX90MjgWNGSuyK5fJlhU
G03IOPvtNMbI3bIMTka1xss8Dx5gkc+xFbDvzuOtDPWp0EgsA115Olw8Q3i+vRi2
eH3ETilPXvwcRsNs6JKbTRBhZgbSAJwu91d4PZZHS6IuOv2rhkrEuny5sgK1Fj+q
82EqgY0Z7UPwu2kt0B/aY7ukSii0PSGUXAv4oAYmVV1zJ5mb67Xr4pJ8yfAY5scb
8Hf5sa8bmrC69BQDY12luU5QHLMtzN3iHh2ZRItyKgVRrNLjxY+Uh7owT8KCRoYj
fQsoLsZuUzzopM40oGXQUtsgaeXTDDMJrY8fDD4sp58KHhRkYTA8I06kNZDnpIIq
S9HELqtQ5iVISRF0a+PSi3DpPTOpC4XIdEESgU7t1exTfJlFHIjN3A2b1Bku143t
L1nXWSHzBnahkKOBxTK3K772BuqZK8mVqaroISK4LtsEh3PIJVY5mVwMC6b3ZNHZ
20LUoeJzy+conae4QMbZiMhbfBSAFBGXKE7EKHxqLror9NR0VId1SUXDhPEcD/PK
tA8CwY4cNBB5fOD5z0eXxFaeNEuWFNga7V98NlJmU9WP00cQ4N/5uOU2fmi5ZCkn
t0LtcTOT9AyEYST+KfMZ+EFnXgw51jeIhHJLkuc94TpeSNXoBIkMHqsu6TSKgQBq
7Tqg10+H64wlQHx0ECgyNvl9rdw7dHnscknq48QZlDev9p/HQjoAw0S7IILzxu3/
F0ND49f0vLRovaAe1Yscwb5HPVvAMiOkNI4CmDyt/BtRJQgPHVp8GnrVCPb9w1IK
HoX87jIvBhN710DSn02okWnE/7qqORdzDEwURWR+Q2LILXhM4zM8FFl7KxjdjdZG
xcy5YLZkF3z7F3WgNtwvPjIupPFYgv1Tf2Pm1Jp6GYgHmKki59Lt8XydA1H7Vk1f
FyA8jmYbAQ81BxxBHmDcjJsUMuxAldkWAPuGs9ROnJFByMe0OygWbOhcagwN4mW5
ZB1GnvEvUfhSx84/FzZLGSG2SvOD7e6foo6NR/WleagIrgb/APTp8gxjOS6Ycase
2C15PAKruDb0r7hqMDmLyqcjSJ4LrFgFzOWQqmqQnlhJ+BTyd4ZM35qHemSxJtNg
ojPdBFfDbHm9x+ELEMAb5P/AJbAFfeh7DW9nGCfLyRKaxAjS/CH+Cgt78nDU2hrA
yna5mC2oCGSqi9lUjHZC/vfqjkMjZf+XjuZ9gzodn/2AnBgFby2FdDnLCnLvOaqL
MfIgq/jcJoS1/6AWJW/RNUmG4agHtPDnVZZt2avZtti56I/icMAeiPvV0gnlagQS
I0i767UM471LcUQDEkyonDRGXNoJbdkVjEfoCDH90qn7RIXOIuq2uGcSQswo3ZrA
8mjqc+K2fAjkkzZIsoektmmaTSmMvTLMMJnFazMGqKjG9sNIoEYp3RNFtuhUpbCB
IqrqFiflwUQX2oydhdp7gORpnHjJqRrzroeaxehvdEHr7dbpj4FC0XcMgs41nhzB
KBzLeUIzKd/LdVANrDpt3qZ3ozKms1Stl+Qfop31+YxnSE3T6XQmNvXLXNObQyMm
2fpos4TxHsh4J3TwacRROLxnbE3uNjLhGoWblF9fbOBXXfDEciCTzRfbcuUgm8jE
X2XOA51FntpEbqve2isI67zPxosI81mx5telfVD022ahSAaDHa0fBsUF/1FCVMtz
5v06PIKD/lucwj/Q9pLndzXOfwdXrcMF/4rL2/htIjwva/rYGWEmO698GbUAdThK
LNDWraJ5Qw4LaZ4dycYPk12WvkhZA9RgxBP0nglPMRruqK0SFLNPDBxRvTHQw2Hj
RzGKWTSeVFaJcyN/6fugA6KYV5XLaUW7YxcgVp2yp3x7Ty87owqgbFGGf+ZyC9PJ
m0sCd6X3avdtM01oT21h+jCSkBykfIJDsDINOZKQl/FF8OFi7Tdmq7xem70eOCTW
uRk1e05bxh3yGTEGr7OdbJlN+q4WcSvYrP9xaJvRYFJn9u6Vczjjl6tnFprU+tNn
Eiv8GhYPmU1pgGxOx5X1WGVvvEQ4wWYCKCxovfPU3bCCNbalMkhS6bmVd4Ab8ZpS
crN0+++EihGIOaIA9wDPMm7cgivJG/p/w6lvx2HR+1Y8lMNq6lD9YPownohRr0pR
PS2rl7aZSglm9J+EvsVlO5RrXDi0Porv2CvQDyQkSlg/mKvw4nNTabCsTay/AwQc
75hkFGT/0O1ElHY7V1Ag2emngsiKd8wFcid9fDyV8JbOMFtSUd6yO/QOlYk0eedQ
z3Dnc7eBYPkhOe8ZQU86luRAZjMrUFjH6XjujP6GxOy0PNyvt4lVvb0GJ3raXtXw
4D01QJ2ddfRTd50QKOcLl+ALMQm4aSrk1yd3GpFs2mKbHO9KtG7XzqeNVmn3n/e0
t3BobIQlENAiGCkEz0e0sQs5M5Lsrb6RjT4f2NqNxv+Vx67HuUc2TFyAtjQoFbuz
Qwp6t/P3MeRyQfByUICUv4Pxo7ar/PLSog28wnFbHBfcayPdMOkbe8eTyT5bfpnB
e8ymA6zec8oD+V+n2SehFrihnsUdZtK8s259dr2bGlviEd2cKvTBlArwycj1lxQn
dRhJ8lZ2hRugX5t2MaWw0rM56zeu6F2PXuBglyd6lxnBcCbcjvLWpS7K1TXFsmY5
eZy3s+RYs+btYD6H+4mmh459g8tOET3pewDnadipjSXsOoKBs/HKIa8pc5SX4JA+
/rCfFL2VJblJ9+BKP3wzC1MT14OnrBRUwRo9DyT0eM9jR0TaJg7oIsURx0KA2ZLi
Tdy41m5ny2J1fJBeYeZKEeervmFaRoMyrjojDL+zcJ++79G4TSl2k2xQQ6C3VdGw
dewMOCob5dJRFT6EBQZmL3eNIZ6lsOB29HxHHOlfXGf32wIbodJbwpa3pd1bxhTe
lqSY0lQsR7bcFtK8b/WmePF6g1B9sq1ls7cs4T+Vwrs7OXF0dmGv7F74Ft2q7cTs
aVNN0g4fajLM/wb3fvAonewv8PE8VQeZJrEVCDV01jDHP+hK/8g2pV+xhPh0aRw1
CgcsvFBnIAYgNq0Cxtt52us+Qce4X4C9+k/+KHEuE0yHLHddespJpMCbazu79Tmt
km2aluVRpA76tPGmGPbFYY6WKMX6mCqH6OLUO0GweBDGUtbS35mzUUYqTMbrYR4W
Gk/L9lWdSs8K9VAAgkvTYMpOGAhIP+3A8WZJeUmxef35CEuxmlZp36M2VPxDGEIW
12Bz9+qJ3/ZBxtnaRVZHkLHiK3wmdaZMHqCEcPHViUjfJIkx4iuV0YZqIMtSaO+7
8pSXgIkzkfqGxVHgc80Rm658Ulwh9BScG54Xb7bLlBJfJ2nRpHYx73c5qObfRAiA
8Lmo9KaY1SXISJsTq/K+x8P9V9Xez+5KRMeyKoQE92K/RdQzsZTocAVmCFAG6Gzf
IhK6kQ3EpO1qBJtwBM6QOsqbLlG+lvlRx0sthwSaHFAZ5cLHnQlt1slb9msM1F2q
f14V00hqTykOaLLU6zm5a+jWfyaTQqsGwjkJk+bV9tZ9uDdimeCTO7qmkprz5PNK
MOqtu+tIn/6YwwRovPcxOKR9nWFcSMmfEhIVZLPBskgYuOkcESD1BKsIMrkAgQi5
pFlXWaKp+FQW1/Yc/RayCcacGcS1yiGU1fnj0riFuD9CTVCGGKY9pCSQK+2z1oJT
/hYb7/JD2H5hTMDTeKowcnGYB+RnvKy5wFLjYz9k9GB/rN7v82r3IXNZfsU7kk/K
NY59Y3ssbAQoJGAB8e3lUOqc70PKNtrw6jV8dFULCIgZYEAIbktMbGwS3yOSxs9w
uiJaQoYOQFkfyESiOOsOrFXL/iJmSu49THWdAPDZpez7b3wlsK4xBubvIEp3g4XR
o4Ou3nTahRMfF03prz3kA7piqY4LXGWujSvcjRe7G2BJPQvCZGGZJ5EJ4SHeLss0
atxUUq/GJ2OpNkZSJtujy3DXStgvejUbRiTFkToCQsPpNgw4/s56iMh/4ftJC5mQ
ONtg09Z96bnj7hb81wtPNmJcGNXyUmvGr/9d00kQ/INRNAUF9wucdiTBDAtcKJ5D
Db3TdzQouXNLBpVos6KjOE3lSTiFvNirb3nEqRQpVsyezyNoXVdX8n/omOwlZKsz
cNqwkcQk0UP60W6AhBSnkexl6e1EfGKoH5aXIj954Rai1oIXytBu6+UOpdwiUgr3
C/+hMe4glW7UKQ0Lf3p594f58XEhSOqzbqGrgO4O2rz0M8jw0jvXZlX78PJSACli
4naS+3SvWlB9u5IJ201l6UIPzrsVnXCPP5a2GVYK27dN860OkGkmxeGCTKC6EYZY
7GRjOjeHxv6MmSr4QHsoBe6WpCE4++SupIjn9f9jVm1DEKIlIB6ceK+XPksOpW9H
64NU6v16ruRLjENbGu0Qq8rfi2OWXOvpM6Yi5iVEjqTEwPTZpaiQFKcck8NuUbjo
p76yl2f0c3+d+wTlMJZU2VkY0xh15bEDBTFZhi17UI5lwcLh5hbPu8RN9WVYauvN
KELufvwZ6t9Ls9LlHfwgJRI8flGEUXgF+IOK8WsuqZFfay2T8BkbDl7ScqUuzE03
iY9qEBB+cGPDLZh3M5qLDU1iuqJIRro6OJ3/oyulene55Sr/xv0vjkFw77jyTxsU
mx8QYkjrI8KrehGMSIpxUxxHsjEOLXHRMy0j38IBI1ZpTSErnMK1aIq8LHapV2tU
cRSdYGpjOJR8sfu7FAM3MOl62qkzMguD3AdZfjkRW7FM98xcbNwZi5dR+WYmDtOW
GhBZtpO5JtbUkSJham4msorNTX00Yh7vG19LJEwPhhkniaJPalmChA5l3FT8MmuK
Wu82iWGdAe0YeI5Mcd38fumBgdkRmVGfHff+t9zHLzHBCFWYOa6YKhLjIOs9acnw
XprqA4ki0MqMFzYuii7S7X0jZ7RU+DMfsCjw/R8mttjM3XUt3uXaqIL3TwdZvzvs
NRfAIcD/B0uBHMDn8RAu/oV6/sJhY5aNEOtIp1LmVe+LWrOpQw6PzQC9/JJdgDbN
Ugw4agafJKq+vGcn7Rq06bUnnJ5/IrqQu7mQ8L15gRHhortQ5CMrGi87OrQUmcFV
bbTqK3PLagg6Lm+tdXWd/uch6EzRyynlkBcRfJOi+nl7tHmmnaAvdb6ODKdGDW4L
000Z+J5fyzTUBFyWFx3kkYFUyPf4qJ29MeclDfKOjdTPLkR47RcQZ0XXzTYann6i
kEfU1J+pngFa4fA7KQOBRBGSGSQMs+6o05jiFxNlPpvx1EoYYCgsAElKomeVpn17
8HLpUIdPW8QyJkbkR/I+lUTMyY6t9pMR/300E9zGvlsgHBur4Q8C4ajLTWgAvTsR
AfLGkHnU2b5UD6jZKxeX6OTpS0bz3jCuTRXXe+ySshPTf2EuTS/8rdGbvgHID6jP
k18XOt4qB/PMN7g3p8Z+JDb27qr9FMKYfMJo5pXTCbHSK5+b0IQXKaB9+o3rd4cX
OUYGXogB04UCLyind+YZNQ8L5+RNSASAULWwq76LmAN1CiPYXeCX8m5Mbi+QRqiP
iFmj9f1cnOlPnEy5TNOssNiLnunwfqLHJr1qcp/b9hc3qlJQwKvN4BG/IMUTQc+D
KJjwPZZO7wtlqavEI34xloRwFUvnBe2PsvHKLSLI1VOok/cBUHn312FPeU6OjmPZ
3WpF5/EQQ4q1YVzN4Bcn75qqY+J75n+XXtqTF4KQPp3QAqKxFUEdGCnt6RmcuvzA
v3Qa9ty/uG3yEvU4Gtg6xCDftN0OlJZDyoco6YDfztwup8W/MsOFOo42zl8bMuBq
eraN15ZM54tYyHVTWb+gVEipG94fo0bUC3HQldCXEzKk1Js3JNpbysb7fl6LWoiO
upt6JfpU/lPe0H5nF263gTlddWtX0bvZqEXQ9unpPwy8uwktd0htSE4hkmGtTaxj
rKIaBbnbhIgY2FvpIZIiESIvq2lZvlbdWakcXcuoYc1zuH3QKzZyQbVujpQmh1EA
FtYhncIVSCptOxq36j6/wIRTmdd1aTZLfUG90om7CtwtBuqV/hco5prpmLueK6Jf
rm5USTL7/zQKKUSQVN5BekK1XnLnhtczOl48U/T2+95C58J5TYyy+1O4JQ62qzV3
iZ/cprYBG10HG6gBZamRPvHjoQvRW7Xk9ODriPmrwc1DfYCWLrIg4kPhLrGQWEw5
o35W6mwFr7ZSXYDp1U9KHpBsvUbegtsiYDE50ZbozeLh7jwwZUkqjROQdeNsBRCJ
VcHbA8AIuI243ipRLCu62arxmi7golLdAC76SVLL9A0wDqFP9pAQeWxYe2tae2P+
bEiHBz7yGuysSnmxftWZ+rUPBNfYeB0y9eaQgKW34XL20RFMyULyPqfqEGU8iUJS
CMfcoxuBcq1w8+mRsm73NBPKt/ZeHnVxFvvH1HvJjELwXjjmdWQvN2ZnzQAkwyTr
ohGrnusi8qesWSWDBQCnhRUYKCLM64RiCAJG0pqztXyRys0Fyg0TfCxie8DC0EBm
32jHRFMrmsXl0Z9DrxfAYXvpeMgK4uPPXJR/Pn2/gsJHrclLnpaqS+o4Djh5SefC
zym/ctD5sB3HAGSfFbKnv2JYpz9xfp+njncNBF+gT1YcrEYKHoD5BjJJ6Rs+r/cF
O1IuKmgCY0iHANma035qppS20aCzfwW2zvFemxT4vUOp6hx9cWN+8N0W1vBzgMX8
OPd2dM0eT5lmriPiAg1J0vL8u/5SLaaCBZPnQKopFyQ2V/7tYbap4qPM5nBtDY5o
5zM3Cp2NzPD8sJCBkRJrUzvvzLkIiSR+BvnOvFJmYtVEPr80+6i90GxDJotWig0s
HwDUn3rrxpa4NFkwTExwkdmadG0TpUyZnQ5/1Ww+wEC+4YIw+9hUV9uLI5rUtaak
iM4XHgDe3VG8LpjsTb70OXc7Vva3C/4svG6jzF22ZRLJfaGOei+1dlVsixcaVbE7
A4micE8rqD5TDkKRaUcxqiJRv9wovgCrOWRB4wK6GMlezGikF1Sdadm/Epq0iwcC
4+ILNIqdaThix+Iuc0eUvUE9vECE8lm+LHpEV53c7c/WIjnCMmWLALIC0oZJF+1J
77Xl+4KbrLgA1KxO1/tfUJm7KEBY9k9WF82yWJe1Q/ezmBLP2qj2VmRG9OHX6Ui7
Dky//4Z3iNO7ODDUSjuaHtqq/NbPcA3vqMqiTwjhdCh8ezgT9HB4PMi67Ja1fBsr
Dp83bB2rVD1xJUseak3qt6bQNzSVrI+tn/Fwl7WfpLsEGUWIdMtDjxhj+9xWf+tg
iUV/Hs80/6ca0eQAsh6UEw5WFYpIjgluCEPAz9u5yAWsSgsU6dMNHcH9EhCKI18A
t9e9l/3oQwfXbFh2T+r4ToGlW6EgMCsJ31CmKc+MNUpAPXTPG0rQkWKcudk+oulr
iFqxedMK/Vcq2zfx5hmZMkRY538miH75I4pz96LwGDLysLXsirc30NgL8jtULEey
fqE0kH0O+soqP+kulKLj3tTSbBxD3m6B/Ora4yuNd3ODonEbrUnxnotQklHm1wiT
NbOfcTXbWbcVyHsqghzYyNUAGjbZL+EAk9L7BRDHxdxgNa6znshtXXabDCdozXuI
bdyYp6oHLhRLDnyHfbRT77uqn6OH6Mr1Yz+GaaxNEShW1/ywmBkFrys6q4sqE+Aq
iR4thLJK5hOiPijV4nWgz74QgMNQ1A3pfytxiPbSnLncT+TpCEv2R+tCVH5V/5oJ
NXcS3zi7HLs3G/vuW6zFBOcZ/L7In7tYtTcPxb7IlkXhNkwNut+DI3MfqYNICQ7b
aBliyHT7nr2s2/ZXhlX5fTE1k/y6JyNbDZg/GmavmfzyfLEsEWFruCPz735SGtDw
96hrbrMDN+MUtXZ8jMHwn0yDUaBsThnrlisQS29p7d5FnaRdPnzGpfVxeaXUxm6Z
UHnFulprJLo1eZGfi7Hjj2/d21XWxWDJWt4QZYkP5bYuYj5gW2XWbpraSJoS56VJ
fEdibGOmtN1q6ez7W8nkfFBoj5eDXacTSZ7oeKOkHVmN5lX2wlZmdL16OyyHqRaz
fdpijoCdmPoWWOs6hK+n/GeOdkVpe5n/wmySMEtubybAiiszKEkg5UExq29yZ/4x
feqYrzla5PihexBvdMf2nEg4ap9FIh3W3bRInB7Wlhto8wDulOAvdYq5zt4YALlw
i5u6EEDFzP2/XAGzaYFGO1HGUUu8qpjR87CLGLT9C4X3XBl32Hl486/hUaS7w0x1
ozrAec8T4ZJ6fJURj9RWu5cloLWf4pzQ/ZL7NftLQ7Abem4zWMvM4ddNM5G/TdmW
JYgX0w/ytNN5OnJyOl+0ktumdJdUwoT6tenGFM63V99RuPQ8o5Bo09nz/depv0gH
qm7EVom1U3gX58DsoHqGuKeRMWyesZNut2E5wEtdEepWgzqKgYuxbwtpUtwP43KL
tNZmZMsQtKzbnX+7KUqNAsOg3wME0EcR/YwiJiA+Wf9x6Y5+4F1M1FMaasSVrLrE
UHwxinedNYsZLtzVCl7jKiSRfxngJ/q2o0VA9g6kjgcvrXTpCkNPPhWKNTZjo1eM
74d7/fKRk6KlVepl95oFEHaoGavI67HNSNE8ylT9Ys017FLjoijQ6BbHVIUgexdv
2W6gYbs6RetvRo52uY2WnwOhY6JYPLGqA44Se8G7iblk5lHaMo8BJH/6EzivS0y8
ft0FPBcyNvl4YUWyaXl/wxaMUHAH+faO+wIj8PuCWTocYZ4EY8/dWFazx6DZirzH
1ELwC0fVSxiA+C0sLF1orFQPFhNdLPo2bdwBrtkdDTWPAbsSn/1wlWfriXJC6n1r
Wb19L+MuSQePpBZE8OsO+piF4TNxJIimh5A2SQ38BS4L6Shv0RlmTqaC9NJ7avaH
tIM05SrvmpzZg6veW+uvdYesJ2QYJLULhc+erUFWz57vhHD7nYesd0LYq5SCFnJV
jtDeXRZtDNq291c/eTlq+OPoxuPryxrn+inVmMdrNJuFqlwB3mbOD34I+5UVPjfZ
cn7XvNZ8d8fen4vh/iiLkXVkISA7jehH1MPzFGlUJaEBsIg+57oykiDmRlByHvQD
fQ5lml4ZoxUOYbPnQmO8m50NcXphpIt4gs9YQYoDeBxRD/38alskNzAgFuM6NazP
hEv/s2x3yR7Un+DrWK3kHHca4hfnnDDgOc1S79RiwXCXwIgTYLPGnkmhxQqr1vVd
CmAEFtEGtzxnWt70BREbPgwRR72MJG+Pq4/8jdmX7gt9eocLQB17Xg/nWerqbm02
8oEy98onICPRz0X63ATqiXbQaHNLaIxCaAXQen+YeZyj3FRz/2PQVUSCGesPiHm+
NfkQXPl42xa0g73iQ0QYQ3QsbC53FcvK85XZAkObojx2/7RQMIwMQyRXFnQQeKJh
1oKw3nHh1sliUxstHV2q1s6l7jrtyVn3bCI4zMLz1XSfErvpgZX5hdam6uNO94nj
hioTznwYqfttlLCINZji8iP7sXHR4Llnyj5DamuhRrCZ9qpmXyvBhA0o/j69cK6z
x/XusbDXC5+iFDOh3Opuuf3qA4XP3BlldpilsSSeBFsytjrhouEhLuV4D5KL/uvS
b1mLYCaaD9IzzIMQv/VR2IzfQ3bJJZZVW5r5sVP+jTEzkAL/vSAlvhl8t3hKvAS6
G5qBlbwrSiSbGjxBFDkGlWfmvh0dDzpFf0j/LvEWdbMGsvyqc9321fQ9wMgYBp4n
7iAP6TVlnmRudr7F039WyF9AlGmwE7rTvOcakicHy2gq+prWQE5IUcgSE/QFzUZh
9+e9I3EHGrvB8ukV68etoC0/7fZU3IrLTDfos0rrAPxcHe4fd3akpXe2tHdZEFm4
leGPEFS9InYtivcPRFLlXfzsNNb5ikfIJWoEJLJhTaK2KccTKmvii6/e2m5X+BmQ
IOl7eEV8lrzkdY437g5+0ShSjuvVvN55HCDUduM1WPBvTs76ZYQMnYZQN7MpMdS0
6SSuDD6Kwg72+D5h06V8XL/l5Ds8lHWBVMcoB3mz4cWdpBEAH3iHq9mmUsxs5P0O
9miDX+hoAB014mZsYQ10wSkadYrzW+zVUPk3XQma0zRTm17jw1mAoL3swF1hXL9Z
bNJZf0eCytJa0NdVeyGiPUHH44wZjMgZfAVmvtdYnjKpuK8Lon2d78/fIqhOOYw6
oCIww9V9n9MMXQHZwoJB3Mgf5BK2h4nNm+fYy4O3BDcjzWDC2GlwLevORfCTjYJ9
Q4HSwGbAXqxcBqzGZ0/u+m+HhEohEzoLSyEqxHc1nG6Nz8BjasiXEIDMjYuGU3AJ
FzTnJNkSt4gQ548hwWnxYZDd9tK8162QvDeA2RfjidmD0nqo9D2Y9Xxai8orvwaE
97NwQsUOhQCZl3yPENqbhFDzbfaXp6nIUJmkC+ntJEV+l6OBTsSXNEUXoCS4Qm+v
CIkNkQ5PZySHcMj4c4ea9gjh8Aab/qWpczy30rzj5t4jrSy5r5ajst72I2wW9B6n
qZwIDXSDcM5GJ2/5EVz8WubpM2kNddYupYWw/4S9+sJiPZO91mjG+9zDjgJlxiNT
qVnrV4d6oL2QP/WOM8yxco0uIPLypfgKxJFGiKWvjALJyiznJwIk+l6eKpWMOJQ3
lOmcLviuzAUQj8mKAGfLLWdPQQgkVvOSrSuDBFkCrAtbCQz4N9O6AV8m04qwl8Oi
NAARzv3teZQ+AfSqPuw91S2PCOX88GvB+brLV6OjrhiFTD9TEW++UD8HNFdp8Z4s
hoLeP2GEpqQbx/J5E+faEtXFIC5+c1m/7P9WzbUU/kZBbKabuPfCipWAliIgh1Mw
rd4icOdmnLnKKjxG3pgv2rsKcHWm+mT3tGy68DjD9bsKPXBOOXNWkQzeuYNk6tR8
YLhKbKOZkpIQqIOdKkVlEwI9AnRUKf+6kAEfsi6qSIUeTsBqyYNTjCiNBlY22bdb
0whZ1+b0mFX1OECB59dLfZld8XXMyf7eMWohIEnhn8qKCl2UM9l5NL1UZpfXaLWD
4ouzSEE5UJql4IgjTM/BqrlC6PBdSp2wvy/2oQRG+EJUqK1EnTQB8uvfO3sRFK/p
51sndkVZjVOa6FWipvZldcZrp8n4pzd+DpNZVG+kQJR5pEUAziGk9LPfC8r751+B
Oxz/UVqAYtI0R7zSNSSVD/BNNUuVqA2haSu8FclvZQBmwP1klE+V4xdbTB+W1n5G
yabF7l9lOemsL+XFxvtcCSsFnfJFqZPQ++CAd2o+io2fsTBVzmMgXb6Hc9qlxjYN
BQed2X6JV4XAG+82VoFGRmLJIFtwkz0erQK6AuC7eJLtHezGhou82N3Gnfq5s1EC
9zeg9GyQGilc1VOhiIDGQc/kRwp3g5vh0EDkJ+GA1q3KIOgUjhnXkWzqjlDEASnJ
/OO1wQPkysSKdZT4pEjTEYRqhk8YORmSZr2fY+vajQXH8Eb2o46/o2vhqjbumSSo
omNF3A4fsHvnbVf/DBqmult81fTuj/YOnX4OW3Zzx0XqHINexp7F3ILhBFKuv5Rm
uaQ1Hn8yosQQHMkavgrJPFDMS8+8sLGmn57SnnSpmP1ssz7P4Z21EsYDHDgE+sKK
AZxMSOSuL8eRYGOc4GcD4t4AlTz6kfLSXOzZEUo3WYQWJwfTEHvGeyNfWj2dnWe3
MLC1DEP00cDdNJgi9FpbgTcjxFqtl1HmR04P0GTQhEqhfuJWBWJ/ImeikUlV0E/n
xVO64fyImeozoUhWOMz4Yo7PPtrjnkLTlBDwccYZoRlliofu+UBM+34VGghrz1Gc
/5mx3PL2J2DBX+ZIzcK2jNlWW9ab6Y2DtxJdt17tUmTUSE3DwDMWVySSIkOTTaaX
VilPbnXdQOSarHtISDE/B5lYmnY1YCYePC3YnuEOpCb2uDtL32HYYKdN/AH83HUV
8riE1dCi3B7aH7ZtunTMg7op4Ug4N9mcXEl+wzC7eimDPKtQV3/d394MEURxAdSJ
D8NLBUb5bpbCCTQ62wE4+ZZPL+XItIx7XKNAZaUQhklPHhSS9dGcnIdbe4ljxis+
TZQrQcRpM9hW+l95qYVL1biaiHkclFX3Yl/wdeaLtRRWsjkCJiAYg2jhEUypw/HC
7oD6klrqVgN92uQHmet8IkmRLBMzU4SUzRvRW3SRJFk5I+l9xnSYP2aa9K05niAj
j2asyP6ZSs4sgcLB78G0tTH7dEq68+kG3SYSNyuB3J6gWkqCVuIk0xiiohvbu9Z8
Tgez/xKFCkofXGLWsYSFVqXDh4iQbTPErRaT1F+gT1K8tJ9Dx5dXezY4zM3B26wq
P6CbmVds5KmyfNlNbnCTcGZA2qhPwq6qvXsfE956iSeFq9RZyuYh2mQzTC6ALIVg
cDl5oyntyiOm3s6cWkC5RkxD7dmnhuob0xSh/ehdZjXTswppyl7iT2DsMmv0rFvW
ogF0k3DUBalmL1g+YIe6B9DfGAqtu36BEdCvi2S/NTaCj2CcMa5JOG08U9ucP8og
LqZvASgU5q2ffzABLIzJVOT3rlXILjte7QEmH21l6A5qFRIZqDI/V82QHILF+fg8
8X3RwMtdGWkrnfflzLLkql/V3Ck/6+x+uGtldmfk1CEGWYJSc4QPtJYXs2MUCrvR
wM6DL0epvu0MO8j9r4GgFyNzd2lMRGjOdvREL/Mv7hXlSuD7KCzFTqQPQ0VYOa+U
3G/whKhh8qd8hGvGOZM26lpyktXQkeiz9iSVbpjVz4vPj0IrTbuMLYtvq6BEld7f
7NH/eBq3JhIJ99bGYFIs8dg6zHhIwq3umkhTTBH0Qp6QzzmRLWKQLOuSvkrIuX84
Wh1v2hvoGaQgoilyat0zgYqL7cko5f65i/ezHtTR2NsaGsibLzn2jKnWKsOo8gNv
0Jm6a5MiUfvbt0g2nve/0hhgd1oNPCqVhn/dQP8dt7/SYi/bk72wMHbFxEwWOjpM
X0tZS46AcEjsNkYkZCj9fMdRu7A0hLp2pe7TrR0MzG7Y+Z0q8tS442Vik86GB8wB
Wbl2DgC1TrgatuzQLGfEBJ50ex08i/rvByeR4fhKFWA/DmB3sf8VJtbuKzW9R8ZI
86ObjhVuFxZ2yvgKpj7dmLJwsVWPOUZ9akNx4DsMZiNSLosHzdC6C+TwOOlMobfZ
bVsV/ga1HulzL4iT+GQeCTmPYI/QmvAcwQQMnHJAOKhAHakRcWt/m0AbsPewAiz5
dHI6CYbygJ0UFADnMxWcWW5Ww/hFra0+PsIR9Ho37lOZaojUkOmXeqgtx0vfr5gS
LVGpIspas/q1gT8GNr4fZwL6GFicwbsEFYCsBrYlim5aC3ultug/u2VQoNYBRaoN
5IYy5YxfLtnMh0fFAt2N8JyN7HGcvjOojoIz1Zper9poqdZIQMGfoyFVh7xchz96
VW067JPWvOOX2LxMEk1df+/2VwF+LsYpNQfYx5kavx9t9dUu6bkJDO+iuclx+lPC
wFyN/T/pAuJcXeRHVyiSRlN1uG/3+CkQy7gQnSwJkEt1tg8CqVyOn07GigrlPHxe
n/diu0wfwl8xw/9NREOTfllHgeUja0JjuWhbaqylgKqDwKCkGnSKO9G/YZhLCvnU
LBFqlVrkG1ZUcJt+XPo3WU5c/ZUPaG4Ann9dVFL6LWHIdnGZBmHm7M5AwgbG25LR
e/JPpyItqM2UdNDhmnr/yhTCwEkywvcFIohQcayfZXTiSv7NmE0lAo0U4395uYnF
YdJ/QKxc/Fqkv02yjyy894uH3ZujixdVp2RvIPYNTL8NJaL1RFzIotrA2NJYDdBf
dfddDDREzn0dFWmoO8CYixojE+c/WURuKyfNTkdJkaMQcr18s6frqf8UtwXO3D1W
DnkUkxzn59d4WEYBYd9dQRw5lWu7lidRHUp4/NilM7uYvQIPG7eiQdNy4NVTv4Ri
hgrco5ls9VbbPkRigEVJ8PkujGEmTj+gX0O9y9R/nTvGCsrL9uo3u/8e4TQ+yKgS
nNLSAD/GUumj6Jy3XjZ5jmJF3iYcOKOd8apUThEDLe9iPGMC3nPtBTLXDDtKd/C0
cn4OW68HhTx4hEmQsLh8CCGU4Q2Aqlg2oqMqOgQrmyVmNFqWq5WHPqqIXt3m5QRv
vr9M+0hjNMdBXSfL/PfroCXD7Vp1rQYEdDPez+AJTfxHnq+UP9lCaYkreSCocA1H
8+1niA4m8ZygcTH4x2W7wlCUEtEsTYrRzmrERZNILyQh2g06NHyMec0mqw02pw2O
KfNhyn01Oc0/8foWL1N8GfnSuXWvk9aKLSgh7OZwrJCv4hOJacKY1MIJsljv+BkR
MbtwNs1hXXYjgobKdblMIRrUQjC7xYmMHgzOuiqymn2q+mefKXT8c9UW1s0drklJ
89VT5FG5tJjH5POcGZqFZvPib6mNfPkcbzkAeOqTfk9emSdm9sfiyUHHMfmGREts
dND9akHLHXrd4A8lHgLv7mUV8ztcGa6Qs0WAJcezodRZFshgyjV97X66R28f3Kus
TGeKiFBm8xiJiKpsab7foOrREbEezXfX38JNXQb2Na26Fc1RfMLlqFG1WVoiXvdi
4j+4kgma1tlMgCkBugvkNaQD4CBid9t19R6WmH9uOcaqGi3x5C6kWk2DHfiAtbP3
0qoEXQ2H+4yMVWB8opQbzK5gH2QcT8YLA7YTGyaQxfqOT7pDGfMBhAq5Ma6kxIF8
QRBxvqeLjQ8ICHN2KeERhFMYEIjbPrqzDnqx5+aILqtLBUSloLrNCFgMjxtuEWvE
P22H2XAgU0vv8NiWHD5MceBn3cIuwrMhKuFNp61U60YBtHdyT1WJJTPuMO4rIPGv
uOzcpQWZMkjf7ftkXBgt1q4Zhum89Brp+mCwv7dByxFI1NAh8BM4q0W2f2bOTzdJ
PvvN6Dxk7hmEyIm86Th6WVxpwcwOPcT0UGwnSoG9u5yU/LLbzQwfKsJl8QZrUbPL
J7meDu4cy/TxuQMITBM6ZW9ZCyANHLU4eXzVz9Ix6yXWjUxzum7ZoNlAtGzVWhv3
7r/SLWpJCUFvXXuZwHUdC73PlrZ4l2f8HSq2mZqui6ML+hVuN8kLJRmplU3ob77K
qlJtq2Z92QVDNxuDsnWBbmZBzMCGOohCR82az6I85oziDvTo0lbr9NEDg8XWQCT2
ynr9ORfXFT0ZA3PSHe6IbGgMfRGTbDuy1qlSsxyCNVZs7GQx0MQHuObLSxBXwCd4
bL1Iz61Swpj1qJx4TSYlF/gQbVTS6D6yf5p/adNnJ3uBxXHSmWvgQ9rvqSj7p+PR
b7310/bzCWe8GXbGp8Nh/4K5DwY3dENFpMOq3GaPxebYnP1WO1JyO6HOliULdog1
W7/1miKTgtGRv9R00UizUxX5JS6kK+MNA2Uv64jZFJ8f/T6hHhgFwtmTgcBJ5YvE
tsCk7uBQ7S5j+r3Eru59LOg+YuUJ4pg1JMRc+UIbopT9qkjYDwetlWfl91rkQE26
8aCLpdfY6kgLSy65WlXrpVx2koNak+Gt/Og0nAoAipp0s4T5ESjyKagxqSMuAoch
bBLUYVz3Zo/7GjY2ZrKbym4EzxtKL0Bq8eYTwD0++pJ4Sp6ymjyGg8AHO7gnG46e
dIDXNbaQmU4UuKLSqdz68X42+6t5BL8jI3WGNfGa3Md2sFK69l0wmpk0fWdv71Bg
YsBgXrj5Imr1OUmv1MniQq9ubnLCETb5ZcKbWRivllxFftM5A4j4ewbqHjKKCn4y
87ysKpzgdGkIBxuMEPWT7O0WXNm7ZfWlFsQnVVjjRVDtkeLEZkyz7bN63g1DpLtO
7Z2vrj6sNvGaaVhhLFxr24QmaJA5IqnWb7jMh0oOVr6W38S4m09Std7hfBoGpkqj
M9BCIs0F9anamodSyrf4Zk7iJZhtvgq69nER1XYM/7lz/Sh3gjpgy0dYULUSr6Tb
oftykdt6JS+A9WFsUbo3Si8PD4kW7FMwCei8hz0jOZR1ZYPaW7p1CEC72eiy/gdg
Yrosm1uK2caPKiCaBN/ECcEqokZsA3vvULSq0enEQV2NmAZLUj+yxTd/uTkYL7fC
xh+GR05y0rwAczdJCH/htxbPWvLjc/1+MjX7WYjUrYD5T3v5Gz19qmNDFv48/C6U
A95o4Wa1AHPQs+PLpmh/K1sstNovqHY0EErU7Lf9oW/sKJ0W+/qC/tGHDYu2Yw9Z
Q/nlkWRiGkZAUJ1ufNXAT+DQeUyiP24HNAn82SrY5NhSTVE3WASLe335r5lDaQ4t
EDhP0oCT2rSftZMla6rAImf6RErMbOhMjIsbpu3uW0Po9OHKGPKNQBCDNrp/v8CU
2S4eYiv4WwiHhnk0tFphHe3wCUvCsGk2QxTP5S4H0y4802n9kqMEtkgQpeE4NmtJ
FpXhSNVgEZqxR4FHE6QOm9xfS/UZrOu3v/gjMae5EJAU2OcUEJH3xwgxAitE7sBW
rSkaUTaJTnumaSMWD/7Xzf7HcTaaJubXAMk+8N9bWEq17ywKFLzT0sRiuFk3HX3/
Xvj7IoONqjqPsReuqZH/V+xUiEXzPzBthw6mkVMd+QbA7skLsHmbnACUUXDBLoiF
hZARmQutaJoEQuxmO8ybgeojlZwua/3en3eFSEcuX92DbBTvB9G2kkFzba6HWF7e
Ky9BPFmlYdHBwrsf8YSI9LywLpUhwyalkGd8Lr5KZm1dz04zKdb2YyOQ9mDJ5mEb
dteBhMt1Cc/pDGB5Uxe5HI0DwYxaGR7sBfCRlZVswmMHGhU+S296N9oLJWoT6D1l
kX55AcbMkviXe73wMBxjkRpbCiB3TpmZAaiXvb75HBfJltJW2ssvHMUhiT7Y/9iC
2I5771lGVDk/Xj1YMqLwWvDAAq8yhsUgT83YdP6p4nrC0VjHE6fgJ6CCbyy6hvtk
3BAvMki3/K2c5hauucwXi5jb9j2l0em0QGRHIx/ZnjV+JCtUaDRz3uZe5zMTDaU+
rARdcUsGrQPH0/YleWfm9evHqkJSfJxh/IwxmoHDINM48AR8U2uTJEEcW+8UaYut
031z+TJSvd82Tj63aGx/sNnMoeZ4yDRMIaSZJj+ySFHHOETGTb05G6hvq3gk4zLz
0oLcifjVVpPAjp1ppvx9LA31MTHs05ehxID0Pqu0FncNjIE3E1EBBRF3VHPtDiXK
g1LiCu/wl+P4S+o64amJR/sn/Izw8XLUVBEdX6mM03y6lFgE6qjWSrDcNa2URmrg
1JmVinj5kGqNeEY1NJafeZ9UEU9mnFg58DXTgKELvMmFXPJyXLNIYlgXBEX4hEIp
8v7FwDavr2AjI1yVjdwrpze4oJGD7yPHJ4u+uZWDZwHspOeGY+0IXQlLKvAtFvuC
rUkfQOTUw20Ho5r+Q+rYCW8nvCzYfWBuYlADxZ7BPu54c9DyRwO2I/5/VKRQDwgp
D65Oa7D0k6c2gZC2RKPtNDmKn5y8Ym6xXJh+O2dSb/s7IiZR+YGGY3eQ3nhuR4jL
KMFYHuYcHuhnBil58Mk8NeKQ6TUFJpjzN+FgiM0cY/PrQS8qQanr6b1CKzw08EfX
ObIgPGcJXO3NJwlxbEdF98KRxMhRiuWtnCsEbFsIIp7cD7U/+e+57Xw8ykuj4tvv
7larvDHgcwgMndMO1y4JKi0OmVjDuJ/it4rfQ183gedqpNoA0w+jE5JbIK8g5Crc
+3BEUlR1usz+dLDWFleo2hLo+vPI6mCx/XAZixQas8OBnxrddk1DAuIADzTsvUTi
PExxXFaIQ3xyFApLp27NoeBVkrIGh8NjqGi277d10mI2pyQzD/WT0/oVW1wdD2WM
I7D54mpdKjel0+O1rraJ1ZNQ1AMM21wzu72EW5TEB7rZrFvNNmlE3DSV9RxNZ822
064upwPP8/BxEetVaTddz4HwsC34fICOA1o/H/OFTOcTV+r8wm7/OJuBdiYUcKCZ
dS+/HQYyJxASonN2DaQ4NaEiEAR9r7mR21SCbwne4X8450NLoU9ZKrE4rovRBjiL
7Gs/5JnkS3jngZmSASda4hkt8c2SVmmkEdc0Ws+ehZuIbfNS6GtVVuXz3NY3NXOT
FrG6XouqDGqK47uA8oaPgSKOnwUDEpl1t4ap1hYYIae23EAIYe2/HDwOUsPJxC0Z
+GmzmbodmAkcSgBjcOCQBfdRE5RuwkGRNqAEmLNmFE3dFU3OfKi/db0f27vXmD/z
C8P2UpXGRYzk+PuaizIUjM+nL0ik5sZyWxyJ/iGYO7+8NLIlBLv5LQyOSw+WnLmQ
4DhIrnHxtH7Hr6S7aVzzRhhXWulD+jBYmQGaOhLbTSTgNKDdL7DFi+pW8/WiMXei
ZB/R1xQVTGHbOnQyiI1lM0vn6czMX/CpVmsZHVlMYe1QUfjiypnMslfNf5IVZ4h8
JRRbc1zhD9W81UTiHiMqkPKgjxULOz4j0/ltRTU9GwmfKeNESU3A979phm9/Os+v
vPP9g4FSHnak4gB8xV745C2ik8fPTobT2RaZEU9KgkxJk0CkTLktGILieh3wsRVB
e4tzzq8eSCtY5T2izxxxPeTzGjYKvQCcnt47n1fLs5vf+t8mHuClWMWB00SlbSW7
FyZlnLhOw5QuOFElG+S06sNXm03sWF1hZ8bxHsTwvOroJsHXd9KiR8/6FsGZ+OMG
owgn9a1OS/SRPCs5iCrPyMYLG+OJUtmHvEFewHu6ZooCfyKfAa3MdE0hoQj1/U4Z
zfSttj0U+vQOnEAf675JgI1LRAhiaKCgQpT1KDkdhogtXzfqHg0gE6vEXjX/ZwdX
wicaV9zvPWpEDKUXfAQEzxujxYev66vWDM7SQ5sm7M3c6M73zF6Am3KovDvCByvq
4wMcqcxf8e9xMuwpGX1+fczibMO4CeugNBg9EcC8Ri/Hdnbdq1Qbi5m2atwe5OSw
eOz30QnMGX80gSHHkyK8s6XpGpO8chPCx5Eham3upqGP5wUvtOX/0FKd1/fmj1ZA
UVuKL3AHnX9iotozJ259A/0Hr46qBr/Y9Iwl1fUhHQdUc03E/hYiSATcwP+mf3l+
5lNTRQnU7OUiFI8yghMRs9zgnqJXY5K0BZdH8pw4N3x78VHLIAXMe9NxXyqoDh+M
yrdwx/9zm03uS0JoR1MPuIkoSVAXxd3t2oLBJSsfxtgygJw5NJxOmOf1VWbwRlf4
1ugDen8RP9HqJ1kjFz/JHS479EeSC6J7fDUUW4+evcIo2HfRMpevWKM2glS9XVw5
cIkrkwGMJ+QK1qzvjQQeifRFEZiFeXbIifoT3ag46PKHs4jVOnd1oKBkncmvNAEs
+gxrQIqQql8m59hv2Z2QPrqgLIk/lQgWu2cM5YPlpAqYvYL1VTqw8Y6cf09WBpGG
8eIQpkEaNFVbN/BX677A1aCZipxBCWGN7hcUY71jspY3w5XJFLhCzrvn+HACd+J+
i1jQ19HphzpXq9QTXTiejryExdww5FEeUMo1EuGaq9XRnAJPriaKfcdY5zVlmNXA
k/UUPk+LYKcnDWUHyDDUIxS/w/79hGjM40Tus/zc72TgfDhwz+320hI6mHGwM/uS
25Xb7y3oasodpCtuFbL0zyyNh3DI25mJFv+wEm4hy9CaxGCnV55+HKG9NGdj0jM5
uVXCcJKeiR2Bllamxc9/ke1Jru58IlIyCNe8zR++d8GB7Hu4B/jbgjTjGwduuBGc
E9L+CGUTc69uK8n9f7p7GPguAc6fx25qa0zJjCyp1UMyGmBdYzVVMvHZ0K1KoRI3
0xs0tZ+/oP59xTRCMDfKeT8JN2KEqR/gIu6d7AXlMwdesOQMKgiJmrw5Fnmzw31h
moBCbuGK/DCIQjFWdlGn+VpT7TV3ibtX9tpyN6NoTH41rpBBRb2U1QtFQRjAvK/0
iqZc4Xt0Gp9AIeQrbXqTbJxG+QK9zHVrgqaMhcVOINdWiVJ86ctkpk08zmr8MVEu
+S9MScN9hTHQ2nRTk5jr+3PV0uL0zMgqBrt0kLXiVqJsVggrQZgeZiwvOw4y7V86
4GhUZx//evpnf0kIaKmIHGWiAyOwOiS0CQCyupadxtkphOUMJoDf173xw2QoGOxC
GAKiwG8o7EvdJY46R8SqktIAaQvtVUJIY+dTfNNK89AzYvV0+s+9zuYYSqOITllv
uIShvF/IkAuKMT1AcELTC7Acb3aC5sOM3Sg88ejba9V1b6d1BN1pA+qTctI9KJ2S
SxQ9/yRI5h1OkR6ZAxEAjwV7DKIroU5+fq/7PzAxn2Atd6SRWa8dJpIbbRK4HQG8
IVQ0F7srcoZpPcMDvaObpGBOFR8J3oNWF+s0PwndLgsd5A4fKMlzOoS4w6BeuPAZ
XQkVN+INpSQi7K+Jz/iibG8vV6QeYafwmYFKOcrxpvXhZx2ti9ObfnEEHkj40KHc
muEvocWJWAfHP/PBxgesBM/aeOIhwRD8R/HkO/teDNur9cVNogDEJzlVX1aa8hEU
7b+K3XhH6smMVa3P3noe2r65bpcKInEWfaNLznv/G+c+UYPo8r98w8kow33HXIdt
lg1d4lVg/bQbDo35Ekalg56umplFC+bGmNVV+mkcRWogIrGwYP3yS0a76+6asXoy
Eb8qQUGbA9rIrC+Ybq0/O3M0uwE8l8lAqWGZJO1dIqJ7xuVyJieNLJ3EA4slzmBN
klrgoW0Hzm/uuMYUB/QEEEBvJNNxYDf5nM8FIa2TfGla8+Ysxe4adCQfH4Hs6M0v
EZ+HDNBM+jy8IoHHFO04x/V6MMnNwM6+GVtg6+s7xJLgUp9ZyHDanr5yduubJTwV
hm/PeZ97yXUxuL6M6DZqARQuZ9xg3qznK2is6eAIiR4I6WPROC2mzkHqguydx2m/
wgXGXb/diUx8LoiO2MT1e4SnWYMxfGxE4Ce04GX431a4SAYFR/ykxv4GgOScblwg
1FaI0OfRlEdwMshi6cLY22NS3dr35HO7c7w37VH5eCQw3aSZfImkUaUbAC8jsXZC
O9PWGXqK4GzSIgqxavn7jaPkxgfhz7Ywvc0/ehiXYhGdiKQHYZynZt4lFlJxSVgL
/YktYP98KEguq0coTrZ9anhIJL+41iILZtMiaWxX7f5a28QiTYHOPJJAbmm51cQD
P5MffpDjE4ueXFu4G1KB8e3scDcm3j5i5Ju+LOpwlewEVaG8ml5UC14/X48rdvK1
IlCBBpYL7MVVdhlNq3I83wWDCPqy0DGLkgysJRqkfqr0ecTx8BG6rxF/l7ZpMCLE
752lABdHGd0GrVxo17nrqroVCj3Sc2ntVgK595TU0s8/o4sMU3EvSB52bYTQP8eH
BkQJGQQYnJx7Y8UJRs9RMumofBlK7Y6lgAhP3KSNT5OkrCfE1uAlIpQoUSQST1ZJ
72KkWnf+yZx1yCHLiqqQ5u9KAHQv/lXFrZTXXJg7b228ckkfSTx4R+/uwLWvGqwi
P/+giHyM8Z59sf5Ftm5cwrl0hM2VwYQ5OR02OzYl/I7nnqGV5rtS/tLjw0bL50Ar
IkQrRWT2w6KL1m3W9Mdp8oWR7JVoMxHjN3UKjNlj7jZMkVkPhdOrY23P17MdJZ0C
Bd4VqUnMSzIlaX2jP8/3YhnWegZJn+nAYOAf9MsWwA1fDOfLMOpuHuY+B7h21W5m
njl5VgfCF13lWMvwIyP2m+FBxR3Kf2NathwqQgQkqLkyu/JDk9YsueaHgzlZTJ+g
K20/W7oOIq5Pg5tjw6AzOdg52crjBsnlsTK8M6gqQ/MPcl6iITpw50UEfDnwHjqF
wq7ugA4mtxsTha1a1hvvUQod78UyTvH9wH2EGA5/UmMl52B4POUbYGrAUlFs055U
jYRz4aIL28gT1T4ISz7cykSQY4+3/pwnlWbQCl910ICNeyGgqGa8eQ4WnGTEdA21
GCAJwBAR9Lt+oi7ybYGFVAwompJizuqxr0759fCA1I+d7JSO2kKEZV4+Epe/Q+RN
RgorASEA7NGz1j/2lBmHSLUn2I8LuVvd7FSCAPJ6bFTIAhxz0bHUXBAr/9JzNO3X
C7FkPKeLSmWAAsFRZzjAsOLVQh/Nqr0j7bymhnKMHUV+zf2e4h8SHneXwEiVP+hY
c4y9dp4C6uXFSi5hbGChA23/9HCFFQj7JZO2VZdHzhPdRM/GOsBJwZcQN18PeyEf
6pr8/YujAJPN97eK7FWKPlY3t+qOTCQr4kla3oeuj/ScDCuzX0av8uGdp/sjRRzi
b582yJi4oS9mUOekpmRPJkZtgf/6rul/2p84iIqhxLm+ANTQXPKbN5ywGdGE7aBN
N4p0e3OqpOxyT17gnV1XlP21j33vMELfkDs49r3VbvE0BjUv/ZRwNYRWlYaiUnzB
Iqcv7rLFB2gLI7O91VpMRJ1qdIVX/C7lX+kdWlp9sVwDQcRgw2pGKBitCq2lgMEh
Z6PsNZwX/1bYpmSzrVfIRRdqFZ6aIgfcVJVzpZ1U3QuXYu5lsFo62HcShqAyVoFY
4oK85KV2PRL/0MpB8QVUnKFJ8W0YBBLO425rzuSXF3mIjaL7WsYikLT7uO0PiveI
En6uEMN3hXvd4d04ilFnEDu3Is0j3faMxrZ1k+8LW4TdDbhEnUmVhWCRuXOGfwMp
xYg6NlPJJI6nb6fLX7MAvT6vcuMsSZIOpkiaLuTEHIL/yeYGgmjCpewuQszdcv/k
pIpko0htaPJVeQvDcOil2qg8+DHKE7YAGXhLu78pKiJTaN8nd8jtt9MNXj8mQXNI
6RhaOXiqVXWa2xonQog7yjWOjlE7u8+Q6zpWZnw4nx+J7dtiedByhz2knU/ViKE8
BXafSlX8+QYr03RzcDhS5QlBhifzvM9YiIEqt5/TykuIJXif/qx5OAABpeE3gIiM
Fz8mHRkWlzj42SDPDVqA5Hzz1vWbpLeBEXCl+XcK+vlIlbre4SvXtRa/3GscxuKH
u6K4ZTSw20l/6JgICnaL8X6uj5xBociPbsPP1WsAOcP1zhTd3f42L1frMds0WWxG
Iw0x85aL3pxhf9lTDQwEP1mlVs4+154rOo+8W95KzIXoiPqzcVo8Kv58Fr/2WPXn
aFu5ZK/jxajbyMYH8LvAhcPmsej8gLmC7+0aBdyTAsrKOmOSYbWFnF128mxRW57l
RplkEGGP9b3jUcbRcJM+o8dLKK2jcZL/xxog0fsWEkbwZoWc18SXIzD9SchW44Zp
hFBcO6Q74BpLfyeqVJ/BGse4ssmDpuL/rEneFV+qqUn1cmxkz1OmIyqqg+70D/qK
UyAKC1rhXa1WELYLMrtsefgJuGiJvnQiAcwYe23EQ3tvcdnS1FVst05zEy1/i0lG
4mzz7asHvhWLaEn73gcTzeT70/WOGUs1zILHKqJRIShFhW98qQDgcuHUK0sbXO38
XEOLfL8DCcJwTj0MxN24RMdzV+UvdQvzL8RT/KgJr0AaGs9loC63ck3Bu5n/iDJd
oMecrwadwLUN2UPpFFYUMsG0rnr5rJNgqXxORPP6gfbV5jeVXE2ClnVGy/ojaPNp
C7KTXJ5ciDdUnZAuaqntR1BuVcSjcewrB+zpApT9H6OYRs53cKib07l8xkEEPp2J
Z3tbAQQRnFhe+A8DPT+4LK+JqTd/FnOWRbofJJF5CSz0ijKA7OTiYQk9wo0ZongH
K1efvWrIariO5zaFnbEqiD5m7yn9TsZcnEUF7ChLIhtinaQotUxyi/o1mGdix8O4
el77CTLWoXweHTcqLx4gioo82+s8jFYjswff0tgvsQm1iBpMHzAdOwSOHo3hjJ+J
Alp+ZOEJR9sHd5R9dWJqzl9oCBDtS6zTJQBTwG6NBtojBgM2JUuRiyAtp8qWlAsl
BbcBb3qqOsTRl2qx2amK66ufxr5XmKYZwQNA14MJLTDrpFpR/tEb9TpiWTBNILHW
OYDVovXL+CzhbzLAn7AzcaQazHDk6Ev2v7CPgGboLwek+riFgwo09E45nvmnNFQz
9XFHzQ8oJkTjEuXExrI3IOXKEhjVDrmQbtY4DqI612ZadRewHGW0tDK73qiQZcsl
4C0JOLHO+SbPfSOVR22vQ4DrSCFPYFG+WOoSWu+AKRMujavI6DA8g8wCda6y2oFU
7yzofbegdAuJXIUcperkSqFmtDm+8U+qapXK/BTKcJjBC6JmnqyBzc9j8JaUS6g8
PDBuYSPtrPjUMu5j6P5RiQsEFOfcr18Xoe9fYf8RMbsn+lmpNjJMuV9C9PkupNCC
ey4+RUGTX7Ndb9m6a50q9AjgfftfJmnxCn18rDMoFlV24XKlYb916yZb3gU4Hdsg
wxhorHhXZVjqb/8xVvWxHd42Tmp5c1h/CjQBbmC/xI2DMX2HjFP3Rh6RjZO4WNnX
bLwYuBXmWLOXhYY+pUVgtZct9oaVlFFpBdyXFF5CpKAUhzERaz2xk74sU6chr6S5
NHf973mbQ3W0Jh9aLpabttFt3lgYAAmWdfs1mMb6cWuWA4WbYMZikVtc4pFE+eHX
nYxAxEv9nsbCkMi1L0I97MdC9Y311OKnumyHe38XwxNwLUX/vANcsZqlh04tEwAm
73b6edFYzNbinlKlX4hrIIcvRcPI4ki40GFR42PZLTK1LctfnFHeIfEa38kQEwE+
wBF4vVneRzGqRhmyWt34h4UVUlTMqvSmTrlUGjVWWATcTxFYuRQ8eoYslkfzfgMX
bDXzltKoKlGu5mkKQ6B1fxlLfdYim2O8fD0d/MSiRqM3mDoaPs+BcKsVl7M5yQP6
b72YYZYR2chpXa2KuWxI6bha9mAFkMD8HCuaNpV0HSLKtkxhIHJB0X2ExspvQj/T
7/NImB9VQRzxgP92Np8GL43hJs1VpwDZib5akIa5VG5nOaIbEynAXaYQ6bNuv2NA
YhOF+4lXCcsTUOg44Yu6tp2W2lbcZxA3EInVayONIGyKDzC6EADXiMtLRlUOt95C
7mDzAuwjZinvaBP0qTJFfDCRDZWw9MqaVlLnjPi35dfz4CxWlq+1jC+Qho1mDU2C
3EbkAj/mzl1E10PMVf6pHRSpYPz/jeWKpDflaj006HZm87LGfppvvGvxDq0IKL+o
+pEaTrri6vKFdrxvl8mbN9JbdeFwSGRBVedXhjMc/FDke0ZgApUs0BThZORIQswb
ytJbwbvVsi0raOtXiK/6wtur8uua5JxC8XdPnJgCBbNWRLi4bjKh0M8xK0TZ9PXf
2ZvM8CQmR6dK8wkVQq1p6ogwr3C3lVACyaialm7GjEUL8850jwmmRZDsl9l8gz+O
jOKKPAZZWftnesdkA0X+TEAPcnB1WxaJ/U75u2pTR1mNxfDvicovXv2QX9EnMENS
gu3zNPD2HQEWYi0ns2Qj2R0+wgIZeD5cPt4UTQgYCYhRzZ50N2jEnBYZIq81UgcG
H+db4SDlleML4Z3t+S0cRTy4A3FNP2NbaO7OI/YCgykVpA+COF92/AQVWpVSPVmP
RlfIm+HwZ345gVKg/auytvFAtT+eaLcxGZUO3mX4M/26WKvIzTkQIWvDHZhytlYX
n1/jKGY2zlgvzROZ/XYCzvqTIL/SYtc+N+FzmQazRqBgvi+0tpnYRcMEYVugwVKj
UXFctgasvmr9T8f/FhQAN1qaa4XrtLtmDck+xum0s+WNQ/8Oe6Y9DrlBDHrofC0Q
abZyhcW0A/bggmg5jQFGVKAjdREjjFBDYAfhLXggzfAqjgf5PCqIO7qfKpXbQxGm
iLiihCsKJYFuOgQfG3hTk5Ho/hULs5UjwGKsQCDKGasVzWHnzxyjH1NpNHsYED5q
1pXuvKUxNWPTltpx0kmrCPXMf1KVh5ski5mXoIquSsNppf20+RH7bvoIe8/XZvfg
D+b4mEZqQF5TP5TxCf6BPlUHaoARSe47PIzRxsfH5zRA+cJ2NsJSANBtfw7bsqej
2l/BTZ3vweWFPG6pc4QtpmWrlWbkphgZAYBPlKwU9Kzm9IB+I/ZzkASxvJ4IwiSX
LNpWAeFRFoUJzdq/NHKgcx47oIUEh2vCfwmTAF1wveLZFq8DMDs5XwFw3zAG4zR6
eZuPdDw8pOew92g2WZK9Sc6IC9JKqRB98oDXjE/jv0gB8m17vU+raQyu406C11II
H/XNJadnOpeLLqQrdRlnyRGiQk8grCSCe7EIXqgnRn/hOau9/G0UVTW3UFhyus3a
6glCS9jtFB4z5I6atuS17ZBzr3RZN27X/LYsx8K6gflgiJM41nVT1GRryGiUu01a
uVyeBZXV3ceidvva9qUkLMKrmJvWxPSHpolvA2CiqXyMkqxQFm7bhka8BkPv/+Qj
JQiRfoUdP9HYbU1FZohDRv22UajUmf9a9ALCEvRFQlntPYESn5mR1xbfJmd2fJtf
+H32zg9B4VYdtNJAPG8hFoAjXwMdZHy6odqJdVf0r6ArFP8qh8jw+6PH3rwClfIK
+eoE5w9YUpjUkAe7oy1kEtsuAY1v+MSmYa5s8UtxXiNbjM/cCucOUPK/B5rl6+gL
rK0kxw33PpQti7u0fCAx9Kl4AyzKmFhY6VMoFZggZu0gpY/sf8IEMOLbTk2DmLOk
anLNcJLq8kAwXlJcG108WraIfg798MKsk6RNTKQLmLjQYCEq/GDQUtQ/4FUqmjgQ
OPKhxQXKMzHLiYrQKfOT35LBtXqm3aSPi+ejfeuWS6fhK7Ci7LDJiFuCQ9L84ohL
DvnpKqxqnl0NNjo88atJguj6j8lhVMJm2zSQ8Jhb1FjSMKclT/tZldXM4PGkPNp9
q0JCwXaSNADB6MUsur2WZwmgy34eu/Qzs9rxGjM4avo0t467iqd6EoFJpu4nsX1H
QouvTMzhUs05eOK+NXESHmTnitRBa77QXL6zw+gpsrwfOauAGWrSfsmIcNuTtaSc
JewX2SdKPfD16AAzQqehLnH8QJTYSnX9ZpZJleVEPBb4YPVP6WiZr3Tq8ihiC6pB
cq8LyTxENwG8ErqcjRQtGl4X41BYIlT9vwsakHq6h7+h7CTIaxV+4Jv4Rstl7dvS
HADx3wlsEdckQCxEukNVn5OSz/khwnhFIKKiSktbmeRCjv5DABn1d1GXWC/ywFjT
zfWHnIYIEuoDPb0lTYimWG+cIPjO8H93RlvNoIaD06+u6scC9dyNoDAivKgYOv5h
B6svaC3RwxHrbVxnHY08HrJHUST1yrknLfcZhzrncEwHcdJf8FQvUreEawkBJ7rJ
1XYVG1xf63rio2FBh7ZXkPi0r06M1wDpCu+XEimJrNaq1IA1qKhNa2ogkW/jxp6B
8NkxYKCCjkvmcSMb8N1oM+G3+WUxhUWkY7V/78vO31EfixpFWc6l9PRDHEk4ePrJ
R6TfJy1ME9sSyzr2ArNNf+HMHQN3bJMNPvA5Vhq5z4SgsViUnllaVadTHijZtp5T
89OwBJUti3/sVVxcvbHe2qDxVP43egM0Aimm4KojhispVZVSt3LXyhBxytGWh59o
Pa8daVCf/4OdKSgSxtm00ekvNEf8Ej7PhQwGDmoFMJmdCus/Sp5adchEEWLKshVK
SrXflxeGsUMLwl5HG6KcFm7KLZ7FXVrvGLXE4KPy4etsFF10VpeV8sevzNIua6PR
2UtIXX798SmrJwcKXEmepoVqXUqIhYu+0+UcpP0CDgnO2QZChpzh9eKA8ZjntVG5
77EDmbZwUarLDf/rMKxTYN4WYmUSV0nzqHP+GtZHkPdGZ/EA3S9swFjCFDkaOBS6
Q0y1sJcA09KAebnhIWD4KDX9Myy5FrnJId4pQlXcaZLVDHRbw3VpTbwGILICrXYd
I3lH+JBNal+3So67VJU5Owyx18OJwWvqVFf30zURAhNqetv+kEHc8Os7kuurmahf
NbMEtfAfNxUkpmRPPwT3qDZQEsbXjB6DDvI7QfbpFYu/bFwV/Ez0OyyThvcWs5EY
qebZR7cfNL79FDiNInFFE9bTQRCrZn+RhJAHE4wUGBQ8xggkGyz91zS4+SS1Fih6
xrfPnSAeer9nSIX8vXtExyNkW3wWFFi/teS0ZXU+Uq8AG60lExr/i4s65mTzzv2m
RtTpS5R19NaOxzK0lWjDPDKe4ANwzrWz0TbHr/36/xXjZaEtTNjZ4qMRX9Z8vVa4
UH+P47llLSzPRvHA2sAbxDshCkRJFnaBtFl4mLM6FsisoT5HB7oKS1mh12FWEuJI
EDXqfuNRw5b0i8YlkoR5rV3+IKHwBEkhpclSi8i7GeLoE3NzqkIpjBd9k2fcKZ3h
TSr6B2AVbKgdy7TcO/2EQjj5YWMY0IvLj7wkzFdyCuUbTlysk3UgMQXWcSdlM+1J
mZYEJ75mwy2GXUnS+GmDlbJT+Wv2AOk0veag5PQo6448+NjeDF+X4UcDJQuPj/bC
NSw7OaeJs1Ux101z+VyD0nQh/yp/eNVAhe/eX4Xd7wufUqixtC7jYGgAJmPKPa9u
mSkbhNtqGkJrZ3UW5+kuFlilqi7mD8X8O49ebMhtMVX2VVCkGMYSbbve+i8rHjPf
2FfDQMP+UBUkUexMgnyfR0WIzSbsbZTrSMBVTQyuKKnaYVzA++LU0kc9lr8erTFD
byQU1HV3E1Fz3p5AKWzRG8EehaNzdvpt6jM1kZQaW9gQk9t78WziZ/kS5raUaoPG
ly1eZtiiaZq/dPk5sCj5GXznjfVB4ei37SUeoZY7oG/vGeIIiQUejXwn3davB7rD
jsH4E5B4oQVAdEyCRatVB2ybfsCddX6TcFZf65+rBofFmv+YXbzq0VhT8vUGW9Jn
9O+25ka+dyXjPhI4RbwAAHMvQe1ppL0+fLseHrpqfW4XemKzmPfEHYY5GvkrFxFn
h9QK/6suykHV+2MwTg6BMCtC4UnPYvQQD3AYv8Zg1yLiVkEkqOQL2o/goRu5D4Ri
/oLtdUxJw0y8x8Vl5v4TJwfkQeqomnK5VbGCZyb9r6E9ELzVET5ebVphujROzEzn
DzputNqcp9mNnTX3FqwQyWpsu00Ylzufbi5BuLDvEeE9xHtshhT5+ci6XTSrEGJN
XPV2gm9gJnwqImbR6yGRk1RSP8pMdh91cBrAER+icv/p/s+fVYZhyhUwkiXFK8RJ
G9tMm+TyAwDatrdLHqnMGNDwLRvM7rcR/NGTzalS4vEnX7bBdcsa1PzL/BFJemhf
wgCGZQl/ajTaBhlREzTDYbJOSLJAkjjvagQkTDxNAj58tvnc/7sa638rqVi32Znh
5Pd4iqvRN8SfqD93Nh8O8J041fyzVgEeaQCbEu6pd0D0dy/8HdTOu4oFO0dNCDdl
KF5n5A9RWHVQTgwg9JU6EfjNmXWFapfbbu28DSp+vJoiUJBzfPBuRB0iSIZhiSUO
tivvxTieBAQ3YuQDH0GoKbkfmxxNvQNdPAk0SJNl5v6i2dh/ZxAib+iRywoVUjsk
7Cy9JfZr/MLkVUR2irRuKBMqb7SMuiLaTlWn+rqvORL5dCOE7Irb4IGPWhFqKMbF
wH9lvZCqO4f0ERx8xf9Po2mfXnfRktZbsx6mBaF3BsT5k8jtsyf1uF7zG31pup2j
YaJrJa6sibXlC0k9sPkg1fkN+d6nmUDHrIhyinvSFN/NtuCSStgDRsGLwLYIeqRV
ayIrBfMEd4ZfTbeOZNVoD/ba1Spjy7MCmg/nPYhIct1Kd1yXz1XrBVIfjCgU/VUa
Gf+qRZ/hsSCDlWRWKDgS30PmIYBYw1Gm/Sgtx1e96mY/bb/508L/dXgiJ5Tea7OX
bXtZs7oYwN2uu4+H/1AJUdN/qblMD8znoAGFE0PrcC4Z6yzd5kHvaTpgzl+Omvwp
onMTvgaM6wqtNsnSWZv0qYHvmQs36nMCXoxGjpg8Q3AQ1xLpe4g5ebYk1fAKN6Z6
sNENUvmgNvBnodOn8MSVMkj9d0fpSRsXxMgoLO+kenXKWM7gmBR06oAY/t6KMS/3
behH+bV1MEs0DFYDiA2Qgt5/BWEGePmzOW3R6//eZ1a92xVqKUKsvEhp/KqGZ8Wa
MHkRBdinRNKk1J8FCZ3KJt1k14pg7woaCwwVeLuCW1ASidrOvmEHM2SYaTWesxQM
jFH/L9A0NvH/5X7zGdCoQ9sym5qv3engAiR6nT5HO+ULiHMr0bdMxhpy3qe0DV7D
S6enZV8ajEgxB5DIcrq9FzNlEWKSJm5U7Nknel+14OmpSy1l7+a4nWnM2pm/6IHe
3gvKoWHlh4YHcDVu1pugfTiGpFrN3p8YfRDEkgMBQ74M7ZrZXqR277Jr/AnEXX4M
BR9y7xoBy+wfFTfFVs7v5RkIZbibw2EtTWy6bDpC0cdUS8qu+hmPXM9iBq0WkZ2y
cxD5mvs101cPH3TRoYBkQhk6i+lWYSRaJjCyNf3Lfd0Kf4ZY5X2yIiH0krf2A504
3+7gJusLD2COfvqx8TbcNgNayZMJFmrfMjvlLHLnqvr+Z0aZyQSvsLhyslUc3HAg
s4BLoJeRCNImNU7y+/oAhDXILm15NSpM6VREN8gZF7g7giF+H+IeY5XsfM3XlJUr
5BLVC0kX4J8BwhW++ZN1HQv/wAiuYM3BXwMMydc64iVOojjK8kOFc9pllo4Oan2i
3hBF8NpBcPfN2mGF449XuMv0YU6vYeFRtDItrBYrnfGhlaw/Uj+0zlChjAAAH0p2
A/2wcz75yJ5yIx7zTOziPLlDhcmX+fDoe3Ge9xoNUjUUmO72j4ZgBRyDXhjBASWb
s8PIuzDCizEcB+rxEOHGdZJpbZ0vCKG1OftLEZRoQveoCqvBbXIsUWdLMDqwjPHK
S/d4qHwg29vuuAOKYAfZX0usq+qjbSwQ64dAsVZ3e/7nM3icGhizjdRD1SDB2Que
JCFlWiB9/ls0KKgSzs9hnD/+hgkU4HSPr8rvAbbN4eJnPIkhIrkx/pYvgIYjJSLU
lf4a5cgNRgtIjnhInTZBbZH4sYxdJE/bGMRN8faAvfY//RSxufsesoqT4X7+H19z
SlUDWATlnd/u9i5aE8PnHQOB2R/6YY0xwOm65vN5hvnW1S9jIwmZDEleeyZ2QeHG
YhI2ssHJGLwz5lM5QwmCU20KHJrcmI8JZJi3U4KZ57NKZZSrgIQqyLsKIAEZ5ZA0
7XzU+qZcCDSDbuBXkfexa4/hUlghm1sVlIW5zBM1C8nYbL3+sBJkh0o4Hcz8LwVq
Va+2D+E5QuFT7eiitPXfjDZ0zC33EmTmLxdPolHlJClHUbXR1AoVlCuNBQpzaK4b
6XWytCZLsb3Ys1XqCa9/70PaH6yCTYWiXCxDs64tmkSHh+qGZbi3193+fR/+NkHR
oqb67v3NdplfaBPjUbbSdxSn5NdslIeG0jEKth6KaEAl9WXTTXEL0exeUyTsNPYY
4j7u52amN88t3+g8oZm3zA==
`pragma protect end_protected
