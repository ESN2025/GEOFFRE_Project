// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
pINHuaH42KsMp+ixc+rzJxJdDNrUkEA8YCdy6iNZF+IaUBiXhaT5MDdos8BFtF3ioS5mCmwDzwkr
fmKSjZcM545V7+D7hCNfthpZ6P6hty8R4JEN0kRCyO6AkWq1+SLc4NMsGXloWQ3HZaLnhoIZyjGc
VnLiE+owXYcgnSeOLiYjYqAAXxq8z33vqpJgw++bzcGu3PrordrMOnf9pHq/7/GrCbw6yRViESqI
rmX9VGP6ulYHci+nrJqa73ZTB4ZiVarqLg7sME5Dyl1dFoig8OOr84/5o2raKq19zhdRkTkhksoZ
1CqqCb19kp7JbHF1MnRjW/vGZjqQLHQgs86SgQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 42448)
qGxVgtFf+BG+wc2+kWGz+Ib6RubvxY0PD3cBRAGHZ3DvlfcCcvq0Xr2hIRcPhKf/scqjTnQzOiu1
NSGxRVKaI+9MNoTO4FBszMnk5FiWJuNE9rgydmv50eLoHtiSBDZw/MOIn6wwQkggKexUIHjucFag
QUReeOBZY3HCajL3NZidPktFfwWHHvpWZfjH3yYngChuBbx2+tjsanVqPglgAGVwlHF7qt3dwl2h
0A4vn6vlaqZ1n3rRXDNjIxzhYFWAe7E5+EToDW9pOJx8oO7sE81h2HqWVoVWaVZrv5akUaxuqUZq
Q9sgUesDeDNaZqJbJhmyngrRLJsDfuBVfqzbzwCeGmY2+vJmtU/23Si+N5re4/Z8v/hmGdO1lj6d
/IHSeNK7LUPhgAEVzwG6t1Jmj3x/quEGppPJEi6QJoq4NBlc5NFX9ox89yTb5Z01yO749pGPrWPZ
/iw54DtWQM1vzY1/VMFwyOZgjAWU9Q0AJTm8i1pmnwspXWlPwD1YLxSGrtWCj0A0dadaUxbzLpKX
zD5uI5Yy6jwFkQ/cZlKxu3YwjXYkV6/jhnH1u+0YpKxz9qW2zRjiJM6m1L2VZMrwdYVnNP21DpAk
DMJnNgynL7EbhtxXlEgmWL0dLDE1Vwt3GVl97aVkGYz4VgR30HhRCYtzk/8Jsw+FnBrb3BDxodEH
IrVXPNT46vHd8pizXQ3AXrsLb3ECfsLRSKC4pujsHdv3Lrky+NlvdJSsUVVElH9ic1q4AB7JSJ4M
nR1cFc1ZrkqzN10AqsP2Ze/YCrQw8HEjpU9gqKECHsSbJbpFknZ5kfa/Nfd+yOpTyVdxtNhSm1cC
JzHdt7jtt75XFkIdNpNM5BtIH70GwIauosE8IXL2kQqNvzb1InMU92xGGihEZa42WkyoRWCjk1JC
pBIf8dySVwBcpq4d+smYijOWcAbFhbPkAc9Yj8Fbw9i0jifMncbwUeYrzRAPjIZwKyi3yLm1dj4s
gE2RfCPH4FYiOaaibXxe9k4R8u2O0tvvPuzeuh/s92+yIMiC54oy46Odg+xJ2rs9ATYXIBBBOoYz
6mJwvJzNYIVCm+Df1J8PZ0bTiTM8Grfn78DL91vAoSSSLyTs7Mmid9NBYy9sOro5sgC5KyWG+Lqg
ArMG7+BXkKb8/h74QDD0NFIcS8Oxw1EW8fSKLonNKepn+Ds8j9nRdA/YFm97sSg8VppbRIIR7aM1
BP9PFFo2VL3O8ckjEhiZiGWSWFNlmLPfO7aESdC1to9050Or0aSbiAoB793v++KzHLhrERDh1b/A
qbNAeaaMP4gK8Wr+DZ/sqzzDfjvych0L+Eo/4b+Qe07HJpW6h8xmEtK6XLqMctQ4kx3E6SNS5Ty6
1fBJMyRtH09JQxiawGlzfvLBaK2/4mW4b4hmg/G2b5v6D82iRfKvYaHSXUDtoaG89WGvEY8YF/0h
bKjDDZ6uk0WML2YIwzOFUC+XTYj5CpxWKcP+owFXCnysVI3qwRe31d7Zj8KyBVvh0RQZNj//nLKw
+pNYFbGy/EDk46ujEGEZiDGwh4u0DTrhPbaTmDAy/f3oFPF7pBTwp2cM93FHP1w818rsI7Ch0auk
KZEJl/jwoiN3PVl5gNwaHHgrmFABmJnHDiR+DvJtQna4qVek8F01RTipYmZUuszIMOnoRkT9OqJy
lsy14dJuZl4SVV3bokInSfY5O7bCynUa0LevBtEWjOUUEHnkvavBQJYxfE92GbBr+/gYdaGB0e2X
BIy/1mUjNEoCrekD4t5duZwFz7GPzSZXtC/IJd1iz4/CdM5nYHgT2zfce/udG+xGNp8yQAH/v8TI
Evknx1nZCLJTux/KKOXVEKkJnWWHtzkJsbZLHVnZWZG05OG1P6fpG//nGofYTuzhs8Ab8PcRMB0x
6tUuj8dT5nmBmpt++A4pS0dW8WVSPEug9uhKRwNhF0S3MYBwf1eeLde5fJMny3fXqTLpwsznoHF2
I8bZrjquuzrBngJDw2cYxYCQb3DSqiNGFugrzdRGJIJs2kQzvwFApH/F/7PaMPGgpBdzwOc3DUGr
6AzF20MfWoITVo1+DXHQQRbIFmXfA0ME9nl8CNrIh2CoieiVM2x1C14paQtValvQVJ9ECuEoYHtn
rWwznLgh1+dAm+ySrBdCDvFAjdxlh/IT2j1BA6LMZnbrrqcOQLTysrj8UVIAs8FGxaHrGlsnwLcR
g+PAumLrYcZ+FkPPL1zeMsRSMJ4scP7o3MZ3Hjpxt/DuH35EPk5JdD4GHpK5O6Y9uzOHbQPCROkT
afC2L+DddFS8QXkkhsl/QOPxp0lFp6mMJmcjafK5aFWzE0uwCOI7I8n4ZJhuVUYYMeZ+axWMZ45p
D0/z/Fx+AtFlalbk0QZ79LfWdBUjFQdnuJ6UTLnzlXyu3oaQQv4KX/o02Oyvgj1P+wve3FomgreY
Y3iV4y35PZEib/d+QcJRsAih42IUjFUWYQnig9p5T3o+K6dv93GRb/DA7YKFcGAUqaYYrMmQ5Y1d
MK+o2/LQ4zwMT3cYr1uYbn9a9LcfajMyqDbxyjqEAcpvJ3X6cVlurc3nzJECGrpcp6TTqUT/LExd
JSwU8qWpu3KHiqdNRXSdqtSa6rJiNYu/Fs25pkqsGQmWXoH+LLKjf7ukCodjhQuOhb6sxR1Y/J+W
ia5C47tUKWCdtkTXWaq0ABOwSPBXR8ww/EzYL9zqMOWQl+Oq9cpofPBPSUInbt4KjRv7ONWnDgmm
oHCB/R3+kwG9tMeCeTcoHnvcbpIgVz9JX8zrFZr6z5XGuS6mM4KDGIaXJqnGZueibnSrrtBT6P6d
qyVbwPbvn+W1QY4RXwBKFVmSjiaGaH896+xtTvBbeB3VSDpF20FkA6dB3CdjGUCcYom5pDoQwmL4
Jx14Coh83ZI3qMjL7X1XXzEOxN0Vko/kZizdodkA897EeH76wFRhdh4PBZTtkv3eLhrDzaxuof1c
m7lB3k5U5+EVerwescpdbFCGhwcKJksBUyVRqZhTWR4q+NRSXXyqEva2rEla7z86pd3h+YDJoTMs
/Acjcm577Mc2Q8JFMwtqeiiAMLugGDhagu1fqcHUmFYWnjpOoRg1eND/9mcO3/ByTRmZ4S61wl8D
30rRJDp95doyxiLHF4YPLluHi3U7Z7cPJ0Qh5kMOYDUhBWw5rEwURwzOCPplW7DaTzKGZU100Umj
6SWxs0Pp99VjpgTJIRK/9L6iy7SyvFhR02NiGs1PXmWNnaC+Adspz9nI3XEySxWULI/9UrzrcUTR
DTyRNDKSQ0SIPw+qlawK5QOz4JNsfv2mPaVfEuUsdS+kpNNLHiyG96gI+RBaFlNi9WGmLg4DQwwf
tYyHl/HLSp8fLC5UUmdXcOyDfq1Bx5brLO3ieTOI6KGG8MBfGNQbVIvOhb0Rr8/G7Jbfg+Q2k1VN
Oy5jz8ap+RRNeZGvnbha+otjCdu8C23tCDiFgOg8iy/W//ofUuqzmXBzt3sJTyXnouj8+V1PPCfV
4F9MtVv/4/MX8/kVSTCraLZpsm1EaFz0c9iGUtgqlGnPsxVl6WmpCQGHvUM4PxQ/PUg0/VLufCdz
9zx97A6uKpGdhBFzLjzKQLNb72cch90gRo6K61k4AMswc/LmgNAzkx12+uj2Zzwwkeo6Hq7c5kxL
LcoAY7JnyXuHZggIlAWw1tiL5GWh9T+5/o4aft27NpYWd81HPYvFI21tub0DTX/YWQmqfssGKPQp
xSbtlCecpbOeiC9zGUT75wLyNIUbKPe7YZAab5ucQBEPzh2B7vaUVrueKe28O7y9AomRE0w5DsjE
hPbSSDUfO57lLXbAZxmOGBAwxI1fwsnPH6zlCTDcbVlD4AyQUTA4IVj4jPEz3uxJKIww/+DN8rht
DzjT3oAaQfQPqMc+DB3q+9ZsLjIN0oDzlSVa18gOBd+4Mqdd0aQ+UPyJ61c66dn2kCxAyg9OvRjF
WhnLMZ7LyoO4EyJ0PSddn4Xgus5D4Nlype2/+/pijSNvmG6q8uFpsq5T16n2JmTjvGp0gzUzYxJz
CcVo/QQ0t7sACOICdfnmqyC46KexGwqOYE0Ij+W3sZr5Xh13jMXJhewsG+Rs5iathKAq6W7ACTi+
M7Qru7erEFaeuPbhkkVfFzHb1y0yTGU6KkiOVI6oHpdIGS3otRj3BVh2NqC3uJgpBF0M72QH4a/p
lfoLEuzCw9wqTIukqY/K88MTi7Bt8N30vhenSCnmamxjFAWvIzTsfjDHjXbdsZ0Xway/jAKP3WZp
xETu5qWkqB7RyZ9xbEZBHiyrQkRFw+J4X7OJw8ivJBG/O2IR3QG4vMGR98H7W0vXuiLaeI+5emrf
MQspUkcKsWHlcCeF4BW1Rfq1ePdwBydK180rHrsxlSpyEnsVOBcTfqBomDX2gqL57KeztGp2dutA
Ga8zbdzE1dcoQHtwhvs+JLV67oBWFLGBz/Sb7144MGHKfTLO4dS3RESpbeAtN1WB8ULlTRjP2laR
Zs5dsKsKZ7eWlVnszqskhMe63qb8WP3+LLck6IOxYjuKx9ufYJM2s9pAD+kn4VXeC/c8JmoMIfM2
cIVMenH0uFQ4eTAEuLgKcGc4F2DIt6xAknyzob040XjrCknKbemCX2irSDOlXmk1I04WiE2uQNpv
ZK95dCpVDS2Rl+k0jcnUZ39rwFi68JTfNe7W9gSpRcuZEVrKGlqW87v8MKrSl6oQEtOY7NnPa2EC
hLYBAYY9g9gZ4sjpqSzJOqD/gjy45SwY75BQ0cUSPhZniPdifZv0qRAKF7ZgXWjluWazxBJqW78A
4HnH8Yv7bIlgzGcvXPjdbReI7OYVNnNRhMdBXp5cYR/H8dRtFlftFl1uo3SsREnlcPJ4s0f94q1z
QVovIN9bb5tEMxk4JbwGDd3uOOjTpnau929Bce0xH3rEWeNxiAeRpN5uGXOoEGvRxyr3PcYAqgyD
ilaRC3rpBnhTh7uwcs3E/A85XFL0ZMZ3pxS3SzycbRGlhdOjLhnH2VcWJNxXk6qDIsWxPDkDmt5C
+3RBwcuoQr5I1VyIWSgZAhyIK9Aks4F+e5CQgj/sDse9qvJnb4Rmq5CW58lAvEwPnLy/vs/5ByyY
wCPFhziNDu5vwwVRC7D3q4W3BtWImLTKcZGlrGwlbrYr2CHX1IJTOf0bWts6Ag5EDPsx7l7ktft5
VnZCOEQQubyYLMI7H4ALBhdaIc2ra6zv0xe7vcpZeEtrbhZ4OX6mnQFf+jsJJkPRIe3b8nQ6GpA+
7UCMOLdW6bECLTgWgpQsOoid17G9QTuWh0vzQxfz5u0bocqhDLY+e1FRl1P9iDXx3/uJ1UZbPqfk
AAQHEpOMi16B/ATlNVTO8CT9eagoIGCLi+xknkIBm/PqqRx0Lr8mJCvj/BDtAEmOV9Fn37/9UUKk
+iu4+SO1jpr6DiUAdeqAVtM/5ph3eYVQknzGwgJ+Kvf7BSducLxd9Eny0gUqQCmzjEcQ3xGaBh0F
OqtiK+ayzIfeabKbXCv/qbxDdLlcjH8UkAF2mbtxWfCR8CnWMrqoETY828/haDOxgknPc0FFUg/j
zZ9wSYD7S56/JPF86D2q+dUNHso8z/p1NkvDiDTRiM2QrXqEOSNJflsGxa9PVx8wtnVbkl4Mew2R
MO6oBJyLUk3YfoQLUNpjw74GuetfRTzLLQ0nCgaC28iGN9k2w9Kvl992C2QCZMEB6WI7YLwFP6V8
I4oPJf6St1fFVGn/67xiaIdA5G5BvVOSUhq2PCHKgV+i7G7f+giyX3bcBIaUN6rK8jOop4C4dXRh
qIZml5G4JtWnRcl+vMn09RcGlqfFxOS3BqHdZmvm0/W6M101VHZo/HgYnqkRjH2tIv1XmfY8/Pq9
SNR+6/Cd4Nh70/IuH96JJQSn99aHkJHDpexPIY8rSWpPZYmYOlDlH+CyDVd+7qMAiIzWCxVeaGze
uEPhwtDG73erK4VzHZUsIJmNmUiJhexR/VBaDRbPp3QN5ebLrOda35bDCd9ICgoMqmDFCL5yN68P
y+koyuwZR430Vw+M71bcNEZKGw6RrPtn8N3k8uqVo6tCvPiOEIWAIHzA8qp+HgxiHzVbnOPuiCc6
G4WZW8VTKcjQOvtbhHOXmOFsnVxpd7JkA8Cc8dq2ggwx4GBYaAQ7G9eH102Xht3ZYgLCafd3b40C
eeXWuOyGz3zjSkyAMIU8e4HZGopXiQHxln+CGob/ldpLs87eIhVeymfh1ahXHs9nQgq6n1jaKMuu
lwSaaD9xPLpfZqg4vmu8//WMdm2qwh/Ol9UgkchgzpqdyLUZMLH31+0VCGaGLuYJODLhBddPnNWA
Oj7cGgh23U8Ol0ql8/7PZ+P5fx/ENRCSdkZnEzEDQhBvpwi/vQEYeIHSAprjSpW2E7qS4bSTazsE
gL7bjTBbxIJIgkRoqKYQ+2H1fNZQSyISl9vKK1NPhOSmwmkhaSARuKBO0gkESGsTDSrvL0cgsaf7
mCYyzWZ48aTweEQOb9UnbFntK2iiTX3y02yMURRMklk35eFa7rcJxTlLhNXRKV/AcwwphwZ2X7u+
G12stxtM9LoAoF+1qdLMpt1p9+spws3Os7RSfuCyRaz07I9BSYALntt5uWLTwXQ6xblS7Ezszfvs
PImrEJ/egbxtfC+mmHcMpffQ9nICP7ebal0kgc2DZhZ8MZdUSrofwbDhShocz1ct3NNjkQWVZG0o
LpnBsnoVnoVz0f9mVrcn4bnzCwlHZvdTAsyRT+bTghoYL6RewKRq3MZOngt47EwUIUJ3cyoTCslo
8Gi7ROXTb87YZZVumwWqz+06njRsxTjitTJtAWZv+szqlXH/v8sKtsBPuDpl8lxJjqRGoVsAfF3x
5Iqd646OiBep45crSsLx38CTUcZjt1dRelxmyJNfuIabHSQFgm63QIkaXvtXnDebyEKYElSIRCJq
HJOQFhlrqDE5jNWXCBG3iJSaNzU3jjGKADksJ1sZBkzA5I2EWWKQkI7BN8gzUz/KTxW0HXRV48LM
b1qAjy/NFCx8vzol4Wt3NZEwvr8W3p/STSqEl/8o+0IHa0thKlOdeYQxuQuyfvk5lT6Gxml170SA
g6poWhVSyUp10HvJPuKG/8gogAnOWWzZ0OgwRuYTLYebIW5ntqY08m4TwysMobPsuz+OqSOpTTWd
rCS6GPyjS81X3St98tBZS92NUFa6nUw+qOHNBMK4dxPI9zRMQxEU/gMyGahs9X0a4iIbszotnqZy
3mO/zzM85gVWrqORLjguNQT57zK0HjEB7/Q0BE6VFx1UhkyFtcNWcfuYc61Vem4AiKfwCJ3+CV8J
6b6WD+1IpFHlEa2LUsN+pijGmMuBIhglreNNv01iTE4/yVXoSQhGfb2816uF+r75LirGOldYCSa9
Nyl6iWing5oPhKW0a5dzCJmJXFPZ8qVwFEj7ReHLQMoiuxgJFxK6vke0WBCdIdiyiUrIwxvG3v3o
WE00KyFW7PHfqPXysvYV19rYGhiUlWg/jF9L9mCGqZ7eyO4bBBOi6IljG6bKzKf/FwEqPzrmAxjm
W+z/fAHTC0gxIKQX8/tCBRD6WfKHxbj4ndkB0pVSYo4bRtjH7KtQ+WNH+fTHD8lj6ggeB69kfd7m
Gdklll8vgmcF8tiSYSqbdETfC5Ch8Bsg7W1eToZqsbqAxRdZV/tg5/dwLeoFMdKayjN0AS27tyTW
BpYqpegFaq5yTOuf7TVlw7GE++jbqiOozAjUjJwPf6wHNB8l/zVA+RgZA/lZmIAPvLxHohuJ7jWD
eXJkoEXJCLIADX6F03F99/fE3utfQy5SdirlZBM2MzihDNjZHLUip4OYKZLzx1SfIvrUqxkWdv0m
w/ARDLLQNgHDxoOglX2k8FKZ+tpa6WIY7UfKvjS6xPUQulb98SWFsTVm7dn145pr8DIGLg04MSeI
Fm3m3d+HIzBxn8cuVRvE1XlGGjpPA83fJmvEC5Jyk5JZesj8+E0vcfB1EJs0VuOoBuTsNaejSchK
doJEt8cqPduMMCg0VWiSccgbp7F1sCPOajkmxlOJbjjz2K0sIjoJTEEWTsnFdFlZB8GRQ8iwr1+s
f3ULs08vLVWr1YX7FOXG0XQ+ngg1UvcG7NXhZWCLou1i8RToO85J1POF49f4mguDMdfG8aYIbpE9
um6Uxl/FdwAgYli989KLj5QhgF9ZQCXO6gmjNFk3eAnjmAxfkWOWOpZ5FMrBXVv9PQ9rF024JuCh
eVZMM9SK8wWxRR7dkwbOX3hJbUBKhqdrXJwgp4xa6+kU4TjlJ5dEU4pD6alqIxunsbizftgl8shV
04W+Vy28lG+7gwpYQSSwG2MpIuPWVRKx9WNQBhp2aW3+AgxgYshzKS5TsGEGjh4vg+2DY3lxWPw0
uuIB2iWZPV7PMrPFwytTcAjwDJnj1+9c5gWNsnDakL/WNXPuUmOiutIMhgrO5XfOIzLIz+DphxiE
DYmjovtWcpFKt/kEsHuPORMJvlosnetL3UJqUJxAYu94ws6hySiqKognKDRDNDlxYQYDEf8+oFAB
7yUBTMbiY264XgkMUZBeYP+6VERtoT1mEDphJYuRpwpBYJ5bG1IaGn43lThbioexuJZjLgT+IIaB
EHowy666TO2biDPQX6IzGPx+0YGttvfyaSoSgr5ZptENVr21smRIfvd+bHp76GYgkQxRWD2LvkVB
RKSAe4K1sUB7MrLV4Pv3vezhLg0lyBpF9mll9xV5a23ERln16bgl9a269OguC+esxYDZbHwY3Mfq
+RLBlGdrWHDCdYzS+sdxgugzrr/tS64dUikSefAKtldvvXmmIige3rwvjix1V/XNwtk2d+LWWQYf
NcVPx8p42BllIoNOKFAAxQcUUjPZ8AIz+PUNWZyp3hMrH6nJmH6DM9/XDF+9SiLZ67msXvnVC9Em
+604mN1GR6WuJAW5sUlNzVfT2Ox319oQ3yPPRd5t35eIOle63tT5AYP1wtxKAKxXtuHmTNd6WzEq
GuC5zjjUA8lX5mb89Q7ZpZfH6dNM7diDTOgWKw/OXBAbGjFEN7/WE1QtDRiCNXU2M3yzjTT54p99
OJPSN9BETE97St524Mh5Z+dptreO7jVuUsTvB7Te0ySEN4OrjkgkIWNNQCgeMPB7OPq5qlzL8/Wy
0fAkJpPJhlskLqqrS63fi/4h0Xpw1mrx48fgHu+z0Yyimhl9b/z7KGnhXk3WMuOb/3QASHsdn4oW
YYoF+z2P53h6RkGIRYBF8Kv4wbqho+8Tmzisgm4Ij6fqXfgVDwyAnI0iUKPK4D5VgwJ61t010u4N
XZzYG4LbSHh3zZlpeFqBdr/Q+7GBGmC+Ad9E3chjpoUEZfQNpLsksHoDfG1K6EsvqKXEIN7T+SZT
cRvauo00l2yyIYZfqFe+ugkx1iRaU/ecNYBSFNxfyXj9jv2ohyA0ona4qRo+IYE4h7NppXr/A4xY
jD6gzD26AEVowzDll5q7sQTwIMbnOCgPSn/BPlHxfgcsqbjiB6e2vgNJ+0CXbWf0Sfdwf+ejv7R9
SXmTaCCJ2ONzr996VO8KcPXIlO1hmEDM8Q0cFYNJXvdGkczYr54izvLqnOrK5HlvSjeJKeNFkLVw
hYIE5jcWceU78MO4oyH0JENyfGcwJQ0UQmSUtikC8E63S3cS8QdFo3f+K6eECm+82jhNIx48Y7BR
475EBEFjVIIdGxnzzu68MPWeMO5eEh3ljD15q3XYzCg9vu0r8BCP6X7GMWFXZ5pRI0nyhBrN3nxb
q2epOEfGj+n+2GbVLmzMjY2szEtcRl48ja4yTNfLAQ8WHp34S0pG031u4biO8JyUfEm+S94bL3FQ
asG+l7T/5tbQnsxVePYcJfuyggd53dgKgv/iYBhWQx7SO1+GZX7KOidD1QWM7J/YLaPrCdz5SzaF
aiTRBKWr6+h+GpTKawhJeDVzFC6e5sQCN6BChO6TlrcJbwTwQWcAw5W0H22KhZKmKzOy3bQSTO8N
zgL4oQXBnUy1xjTJSv0h/PT8z6dRQUHzLBcGLoqJUhMJkqf94Y7navvDZF2zHLSHBuJCfSoHefVb
Zg1cnR0+fg3KyQ3Ik81oXrQo12e22rZUGg54UkdVG/VMPR8OQaDzBlCd+n+jAam1QjUQaaGdb41B
P6u1bOtJ2pjrxmscATknjcD/ioiIaT23BirVLdOIdPkWh2rFFUa87b9tgoVPyCxGH18yjzJT7vKA
iaYsMZlXi07YEibidx46iUFBv2KHVIZ2SQ+yjBeVADuDEE2R59Ukfpz1RtY97EEiXksKFXQ3qaOq
s6xN2NKjqX//nXP2uXVOy08GQpBzH2R1vXQtp1STsJuekXG5DpRiKpj8bwesGjVOE5rVK9Hk4yK8
Quf9gWjNm3q9V1ese0Qhl3er52irgYy0NymilMRSrqLevS9OITuDvgYfUWKJsCf/0fVy9Bp8BNYd
AMCRGFTeScI0fBt4R31FZwr1ydgcMUXKnI5xEA4o2edMEIn+owN0YJHELNwFyceYF+3BAIdI4bJ3
eUNgEEfzW2hhcaBzPpNEbr6J7rYe/KeLlwiR9dH+VnYChFZ925TLARMDQogDqNGfxBYtlY629zFa
GGYpwKzYdgSZksSYcxwbUAWE5phBbj/w6abxw9/ImMZhxbwVky5P6G14/OZukBo23NMKwOY8Z6vO
D5wZwLCRepOjRqAWlWngzyqfmWJyZT471yOk1gBx3onDUDzR1hUgx7/rmXQf59jvO0QmM6qIO30o
biA0j5V0unHVdAqDaP8XS8Lz9t0ri588uPCP4YYRPIt00gosv1h4qoUMtlOpQnfbv3xkWhFgAmEK
7bR6wlm6zgG6/H8/IR6QBdFmMAe6jxpizkfWO9cGc9cAU2wOaqYoyIdbva9eZ8r/QDNExZ3foavk
B+Jt0dKKjdnTtTDfFQRRNiBZDW+ZQIOThoKpEOmpdcxB2sUd5wZA7/DRUMCXY63tlrO7m6lAfSot
sVv6E6dByoxeg6cXfYRSjmtwZxGjqYpUSNOA06gMKFdZag+qHvcWjFnxvXL9U9NCE80jVVButjbQ
Qe4M+sKhS7w9GHkN7P/f/f5RJWFirno9TyMaOXHu/cNOfvDDSjfqG7G7npmW0UaP3b4N+fYF3cSe
o+DdS/+P7QQTeD76VV3LY2iyXM4CmUWhSh56imVoST+kV83TotUBs+5l2Tbiw+fSVTHtISK4oQlK
XHs9YaqtqpBGUAt6N9nC2+dNIcAP5L50VQ/Y7nTny3d6rY7Jtub7x0UKr6GtEPizZFvlD5x57JRo
zJzII0BDAbTG9RsFd3Rldao9ffBxP5xREPkKwINAoQSEoiJ3ZkPPxvLbJlfW60KwkiqID7SFdUmN
HnfHG0B+eqx16vGqsdid42b5NI59y/cPYb3SUxtF5OfuKIzGGQj63FEARW9iieEJiW/g8xCndUHp
gRV5l5z4vLGXQlMvO5iPYaY7Hhjk9TqERbo6jcuecK4aT/s/03unGma89xzrMtEG42pObnYPusKq
U4M0NHLTogR/1Q8PB93MENsHXReubNaMAfAgO4CUgnkEi5ewzYB5XQWgDM9aIZbQODhagkYyDc/Y
VhAM4lJW/1Hw8WlztMivH+Fu2QZ6H3M8/MH4XZEOMEForUqE+8AzmzCzzngitpvw+AdoYKJ8k/PC
qbrrovFlPxNrk9DSszTyFVymGz8CfTb6e0XVUu9mZgRDm/JXtwp2DcpI4OjDHiV7KYPCah9d2B+1
7zRL7IvFMqYYcmXtVjXsPLM25As7zlfPhD4a55H0XSqPyEMAEVpK3C8OIuqUOBtdAqM2dxKgH4oV
cxTfmZRghnmXDjTqQMclPjxM1MfhNuCjZuPULw395+anXBJ7boC1GyEswnfl19gQxYYtezCNjgtJ
lOnAoXKHZTDTzPklL5aKn3FNGG1F4Fl0ucL/3Vc9U7Pfhm+vI1HUJW8Yx00NoGIuVxi/5UuJml3h
Ak0AWvheLtjE1YebRWB+kLlk66tW5AyGCMG2lZQshRpEJLXnJAEJD5TkYE52F+h4ptc73y8TbDdW
BHGwKltZCL46rmGHYrUIC8h0pzy2mHXDfvH5ZH9TVVLFKz1/XJDfmol4npm2KGGUe1XrayT0BxNO
iwn3HxVq+UPhdem74Ttw9Ay9o5IP9t6pii+TwrazFeJZfR4VJeWLiiQnOMqYkGWseOUxi5nvk0+x
RDB6yxzUkqEIiEPCZTNAJlOtj2Svaybw7H+2CArJo7dEBkGmq5JWISjomqU5W3R7HUOybM6vEXq4
U4Q+D+bSQdzf0guVs7MZVZgdYmCvKXZni1Kb9aGqq7ZqKyWT2o8Hat8T+8IdquoihXMpdI5x9LYr
HMmLW+3A9OL/w1Dx1QZyqBetxsSBZhqSOfE0nIdMnD3iqaXiTZE/KizbIllvMRQq+AChCS+K1ZOz
u1Y1U15s+9PAAjoLYbbDi6i5+EWy5YRPd8SrxA6cVl9Frxtbujnywz3b04GASuXiWZjCuJgAZj6P
5deU1ydmgIUhMEIzsGxNfDrvllp794j6xnG8BexhslD1v8yp74snAzD7SaRerlmf84ssPRK/Ebrb
owbG6R+dSfU4aEFD1kNBLEDwcV1cCbvvWFkLrlmH578HZLO1rt7mI5ivyYNU/lsbEWonrFdtSMG7
gqv9ajNycArlziAw/nqPKKn+48ILyEXC+JRvRuCF3ag0ELcjY6fnqGI4dSj8xEjSWgnCPVFDYpR7
2J7eKXIswvd1gpS3aW0kpM+Hv+Wrd1OrI47OkMN3BkSJTdMHKgkXvOFnejvksZE3gX0UrPrsQPoU
2DbM6gELLpIF5QIMNVRWm0N6XBt0MvilM53PBtDW9D9SEnKbZDA4R3GSQvDxT9nanfPf5Uu7YJ6f
cu4CNG484/4Jomo2sgFj/IG3Y8D4fP+LIV5mfKYkbaWptbzhIeXefzLbobSe6QsB2bVHprFlBY8W
JRj9kRaer6QyNG6T7sJlz+eouzvB5WMbLadEliBbo++7xjfDwmyT2SZ5hL55Cxrd8/WvSKT/k9Sh
Q6jLaBitLA+lX6jLrQb2uEq3Ul2OxnA1+WnwMKVhq68uEwoyxzgrvJkpq1p91czfVEE7sQp8hOF/
bz4RVUHVomcnb8KkvC5q1aEWx3DUVB0uTd6gY8G1jM2yzNDTFC2XpvaNilkfzxA1Xud9StMgpKT/
PO0aIHQduVgaQeMY59f7nCecEwG5sHlOMN0omekz1fgK60fSVipmpaVEvDiKdIi2OyAWMqixcg6R
5T381EFCO4ppN6HpFreiDGPbi9TjdG/ZHsZsHURoJldcidUZCNrEjP0iCgncR2jzqTK222KGrv9Z
4Ag6SRDRSzZgksVFKaKYwIos83Z6BpBM4HXxYHd17X3a/rH82Yuk73CKO5KI0qWULv197icAJVzj
ISNu3Uml8o8BPWB+KnPNvpVKRfwQw4ewugqyZVnEdqk41DArmoGjNEA/Dp8tcp3HiV+bcMByLbQ9
g+RmFsg4/rorkfsJJ1RnJSJr9ssHRYkaGpVePSPsWI4rR2Xit3YP4frUx8LxN3+mLteOLAgpCSQj
oDMTgcwsUy0I6eWOd++JfT+AMUC09113rF+Yqlo1j9NX2CMTectcRz6mt9FDIuQw5/5Ri8GJqtUm
XszS9eDPFeg0ZRbvut4gqsUbAa9hbRDAeQMtK8q6i9uNN3Hup2UUJSJ/Yw9cyX0jISG/tw6ZL/vx
YoT0UfMRDdFfHxE/4AJaohYTbGz+CvdxiOQ+sLuxfRmyLz//3Y+/ZLXNakVm+dNOurgm01M7Piwb
JpiMqCGwlgCwNf6BZPmGcKGMArM2KUGHp3G0avlP+95gGKwnJEzjxhxfuzvZBelUIlKzTLChSqZ1
QfxDAS5eTpRH1LJ/+SByLchTe1MiK1y1Ssqz7lA6+fU4qntUrfJZpUW/7k3xqo5DlmOl/KQM8ee3
7c3wrQ3u0rg/H8snjcSNjSM5ti6Ue1z1xPrET44Abkrq/3bwBUY3lntwdjW6aW/eugjpnf+T/kBY
IM8gz97Ht60DiVlG19ZwgUrfoP4PF72k+aiVwid78C0vbjwalA+pEzRVA944U5WDCwiR7dCsUo/m
lAGKHcenG5kh9oZvxdHxNorVB70UtKKTHCbUHudko60+n/GEP004hIQqBfqBFerHarteEV/414kd
J+siKrt7t7dzm87hnR/S2E0h1uKTE/MbDU9KFr82YAptQjItyjze5g+UEWcn7IAoek8sm4UlqxW7
EuBk8zHwLmAyqRKAZerX4oMwvB0j3BUdaXC31tT8jIfs49bynhrC1A6hL0gckLMlnIrZUPmBJ+BI
Z7pmtsBLE839Fg1WGq8QOVZqL7kMkzXi+NWFhXCAN36xZ49WXtNoreHlD/IIBXPwt/KftaHeKzEG
v+20O8gVAoGgM6EnWQL1hz1ekoXvLVNcB91jxONOLOw9rlt+bdCxuCFhOFwhVmcUgDNypW7yOnE7
BnrB17mj5DYc6Cb2YKKMf/CV+mQYwisOncTGAQSyMTOSWy48C1+jnIiLfE9RIOgRTghiim0wadeZ
Fg5Rg60bjUm6I4i4lbj5X57Cy25HwvtuaV82FUPinIz8MlM+BBmLhbJ54pFwwmTqxcLm6BR8PztC
r1TK1gnurZX0UVISnvcI9fGc86dKArb6FuqQGs+TYtTvXEiEQGrTDR+SUAkt8l3lkT+PRiTJfrEK
W+4vIQOvt1PB+DhLOFDD5DI6j5eY/O+lwJxKTljAOffnERyyAvMMloWtRwyizLXZ424cXXcR5llf
knmOyEZK6iF6rdcLF2VV9Wgm5aViH45LPEHqb6EjCyY6zP9SSF7rnDwybc3q2ho4OOt03VuW+iov
dIyBTg1NiPEGQv9BXmw1aRbhDaF2tIKRXL5+Q8TXcm37QC0/OLiH351lUFwlQxbT8cHoo1TLAHIs
iPL6M5DsJL6x3hFRGwlKH4UVuSS8W/4qWChRAD0lVblG/IA8c7pM3CDgzBOjKbBz8IQ3JMCTuV+4
QVI+Cis+1pYidFva1xz+mMFnHQztAquQTtdhSgvY9LAkScigVqxCjBuH0cQVAUK4dRojQamN9Ocb
90s7HU6TuExUxvHRjEpSmjJxyKN0zwWcNNP4LVeu7WDwIKvYo0kfwqUsqRMZNHHToHmCWW9SPS/2
I669cc00r+KgttpNREcLBlQI04C9cQ3Xj2WHBj7XgXLmL950JMSzRT2Fz7UQsRUG/f3WAiZwxVbe
cRpJyxWyprDxER8Wf7OPxkfve72vvp3Cr0Fj38H+wvst4SfUt0bwxb1/Q36n4hMJZuL6Sx/tW3DL
xe75QAuxk6QtAcP/6ov0EG8plnh8GQ3MIIEykGJ46NU0rVeMEdksRNuSHD5f2oB6CI8WAueAXuDN
ayEN/hNLRdNScRswRckLNUowdKVnbfXd2kypfxhdW0HctwjBJSf6o322lWClHinasYeFqHJ9+b10
6YJa8qO1EL3/ozNQPiokIaFH4O0oCLLXpPkLv1ZGpJ6h4HDzD+vmE1t2esrYBHF6UQ+dlISHF3D1
6zPqK4PhgYH30KZtgsTA4Y5cVY8NORYq4Zgk6ccQd/IuOSQvlwYGW2GzHkDvqcTWkLyYZIQCmv02
I9JT8Rl/sEoIp9+/LgyqwpQAbtmldI5NFMDs2tpAzaVxuj8WhrmDylVGfvfR5n2E35QiGzPK0bLy
9hzMlLnxA3unl8/y2Y77O83GtzQjXIWc+0Mbbzk8pXtN2xrgRXsfSDoBp3R039438rz+q2EsJXxB
x6HcxY5E1cXIAbPWw8ZW+fRd1OJ5K6MSfGI8bh0R/+Ia3YM4Jt6Lqfxj9WaFltAFVbBpbjU5sCgM
m8Cq9Qw7cMpPWK5CFHvERBe4ysPu+yMHXs8ylA+7U4hPW2PnfDjOOjulLu3HYkirsKNyFNGXgiR4
ZkG0D4MsWF6KxUfAuV4oaqr8uMumE6/hBBCrFrbZwa9fwJSvWbJZpNGW+aBDfAo1ORMD+0noHL/p
Wpls0uHox9KSOyKOt6TCqdvITF54jxmQSclMI6fcRr5o9uAC2hyc4BQAcvFvgQ+gLqxOXNqky/Rd
JrsXRWRWRSKYWZj6TjndFz0GtcTNAZ2D6NlP7sbL00VaizjBLIqTqY+DS836c/vo9/aRk+aep7yS
qyPjt1wnRWVn/8eWBGfMsg07WncyIT5GH7H2duayamwxchJkCZPPAdJ1zDhAg47vu1VIi5eh2V2H
yssr6tIqLS/qhREnrMVzpAUno762V44FOHquYra8x7x14LMKS3GBg0I2Q9714Us0VExyVvjHPDGa
o3xFtzm/WhiPcFfR4onPEicuVs7b37Uk8gyDAmpopZnTQL1IWnc+D9i7BvXVShe4qlwlRy92ErpS
REQ6q6CB2SG9KhUrPQmFCUMGtdisQBsxmjhhxJ1SarUSWQUo6dZMqGAMaArlZ7IWEjxXG6FkXQ70
sVBenfBxVhXplODHcnvZDqqyCCBksd6dzG0z2SjJna9QETSMyF4sWwsp+gkwzKahqttt37ElAq4m
YhAKNkkV5aHpptHrdiy5yyMo5tFgddt2+jEk0dMMRZBC6QtYg6c1hf4iJngI7MkwdvDJiGJUJViD
D8wgMNnmfwnbLzu2+e+YU6m2LHyXlSkTbJ8TQEhcplF5k3P8U3dlU3FOnAnhGaG/KoXTe1qDogOL
/bHFnP/x5cs1mFjju6HHnYoq1bpkrsp4tXTG6015eC7FKxJ3IBYv4YHJ5sC5oMQXazk9m77Krcz1
gBarggJIUy5zV4aM1RKoGHs091miq38Q1FJ5MaFebGWIuXi+haRwYAd9UffSWgXnnqarGR/38M0S
zgJUghiERJvWRGRI1amCP2VHxyj6Gx6oIbS/GezLkmX7b0VCV9nN8M+jdE5cn2BWNmA/2nXkaOCn
sS40ll9gwtFf1N5e+xrtZieesrXfQUx/KJxHCsPTyfzhYgXIwQob78J5kWRH0/F0gfcM/396YNCP
EgMS1/u87UN1/Rsuux9oUSxA9Sxc+30O86YhBvOD3gyfu++AWjwdH+8hp/rhN3n2sR0mvHeYKyjn
4hCI2qpcjJS8cZWvsHN20mqQhGSQ1Gwvt1VEqEwlLPQu1Sh+umjxGXcwSoOh+ky6RKZ3JnO6PLB/
ogQzVfNmQ7eOo2rQuTg/P63ELwOA1mkviAd3uPeLYA1iEXJcqOGj+YYc4JNQWW/lQ1pivg4MpMup
AkBIkkEcAAgpAi+pwj9G1wDWflrX74q0H4wDNOUHd+HrMkfzkYfeqr7Bj0qQ2b43oof9HqGLTB65
lB9sk0LKO4YrDpL1zDJW3vLgJ384Qpoc1/EvD2SE9e/Jd+EURm7L0AEjWeB1FQ7RWL4hzhu3Sei+
aVtjfolJ7JJIrm3OlTVlLdjppQFXNdHJkO1KZmCv6L6On1pa0Y2jJxgonAqPA+PVnmg68Zy6//7O
77Xg12iMlx4v3l8Nt7YltfGc273yBFD/o3O7bHS2gYeemKt0EeZtV5icHNPOxXg67xNE5ceX3pij
wJMpF927872/tftbiHKzHSiCCDlwnjA3E+iPCRp7IAmWm1W2K3VQ8AVqL0Ph0cSyn2oIemR5tqPx
1f31w5TvQaFRjibKxSoI7C2kfa4pnnz3R6HhOCiVsaFJ8Irs4OvDHm7mSochXfurUflEI/iKaY8s
b2MM9uuHMAzMvW+YZknlB6lrckXNUWRPhoSYkaSBe5QKtzj7rlDYZaYm5QYLxglLDzJfZbmT8nr6
rMIEqatESy3nH5y5XHC1CZVMgJXlF2QjgzDqzszmGrfZzTlsHfVlwa2YAmyqfT4diN13HsmvL4Y7
l9wh2puKIp+fvu1N36jS6LIRDTBMNueFegBqvsZTLx2BMdAXzlT0UhhiKIUtX5AHzhKnKenvu8+a
DUTkYn39UQhkEK8LVuAD2+5Rd4Z8jqHi5DqVq+Rcb8jLvarQ/dSN53Qa65bw/IT/jMUeGqbHx+DH
hHnKOYGUP9YLkfU/Y7Cl/Oqp7bfggb+U3Mf1UnP3Idrfzot555zCFJOMP0iTV/cViFAL/fqyi6kL
gh6Wu9k8JpQn4VVc3H4L57YWL3ZFfOX5NJt6caDfll/PnWY5ArjmAO5J5oSVgwQFMyWutZnRWLGe
KzlURX+LVPtEX8BzouyyPetScGRg0guxVW6CqRV4J3zH1R6Vhgqs+7NtSIbxs23jpXENjZxoibK2
z/hdjnpo4mSzeNO7AyPKU54Hme9P9oO9as1HJTTeIvpZ+TMImCJw3VKYt9hYnzp0nK3GyPfl8S5R
v4iefZho0f1FHiXPWJhJLBSlSJmiptL4+Wa4OFYi5HN0Psx4WJStIj3bhWiPx6Ug7xaoIzOJVtEt
dQdmDdavBc+5t/6+iI6O79iRWR4iXE3iTIND4+bFpDa1vsTuwzjQwNZc2fQqf/shuZLVHjF/2Q57
4T/F7QwGGN2dPCm/4tJZ8XYOSrWYxDLSb/ExcWsT6+5sMrG/kKou6BhYVW0ZB/kiBqER8rSkzoaE
V5CA0eAyrZkANR58pXJVA7OmOyKDmJIgxx4oDm9glY+D4vEChZ1CoVOLQNfRMX3SapmPIVcYTMYR
HILAiV8pMWBxL5GQllchThC9UhgW7MxTTXaDAiMnePXA/cupkQxuOUIhwRoKxpEUylJ7Jv5Y1S3L
BsXY/9uHmLYYyABtWD8/f+iql4HnjdZOt2PfRbNSR9JZ2Hn+u+0wiiKK8nRsMixOG3HfRxkHza7n
C28faz+pJg1Bw0jfMeLN5MA+TFEmIyKyS5uNGtIUIw0e3mtup5i4PBVmaUVYeoyPZhsisX2XPX2U
1xoSyYDaAv+uuJZFdRg2gz8YEVA+aCPyztwydp+saxl86PJsb+bWj4KPK1W5DhzufDkp2D2gGrh1
mrxFEh+xbGKqrYCwpU3Uo2EuO8hg0Zo09HLa4hb6/lrgjKBUJDtGcPSAdSG2ot2usdSN93XlAsJq
Q8z1mgTb9tK3uH1fwbykf9AW0do4QKiuwVDtLznFKb2ZN6xezoI5WJ87ytSZCudXCtpCmruK1tgv
kDXOUt6heRIh7GycHP3vgzlCpUyAsY116M5rPpWq8lOFB6fxD0YtlBGGUpc2g7+zob/9K79PgbZx
rJJZoEQyngYkK98KvK7m7+G+L8wnHYZr0YOU5tnTKrTPvVTRyAxYak5ipxZz6jvzqNxJN7UNJFUh
3Mdw24BSw7zjaNq+t+nvxRTJt4KU8TuzHiYZeUPeu1p5Zjzfvyq05xL2yd0WxD4qBQLKQ4aG7bmI
xSmaAVyRyJE1jK4T1R7Im8+mzn1zvoeEmqtIlhqQk6FQnI3w/fueNvZxZXrJIZApLgre7a1LbKui
MLDc2lYBNoeqkzb2PjcGix0nbcHj8FUpQIZnCV1QYv1X/Odfyrb5DLC5ZKvekvm/zrwN+yIP003T
LjbXFL4x9xCQGFiUTNYtSzF1EeytHRzhM7A6z0BXP4lSJuAFl3hPgFfFWv351mDpv5C1KZy0SBrs
/x0f/CiosS6hQH31R/hice+C8+oMx08VkTGAtHw5TEdEfEN/qhn+Q2iY6RfoGIkffJPfko7EEzw4
Dtb9GNoBj5JjXyhz9Vb7pRMwOlEx9VvKhtOqkGmlvE9pfPyI73rJpx1pY+q1XbhWJgW5bZZGsQxq
990OF6Z7uQ4jpZL4wSqHhYThyHW0bpIyzm8jv50K1HUep2ERR0Tw605MsTppSBmSqnYbB4Kvk9NL
22lsArOhKRAEEnP5jm9N/Xj+4CY3Ez+bDmmH9Hpzz+x6PQguW/j40A5BIa38sfzMH1YYS+Ffgeu0
4LMUL51NO84PKGzO+CqR0IPMBIQ8dGsEM/Mqjl6ZmZ5x07Ib1xHL/wZiNcq0+EaosN5G5IAHhC0l
qlkQLBVuMMEapvt2Hz/UsJgZw6FugPlSokoUjo6gw5xLVLR08R10fFHFMbCp+QsB8FI7c4qdKcEZ
E249PUSYE4W7Mo9L9lG+QzN9sHy2/B/JOUTlrRBWFQ4/OFYOZuIEV7NbnuDNWOwlKEX1fQQuTjhW
3afjatn6vJdd7zazfdA3JXzwmOE98gq7V2Bz+JDC8Ly93wL4WiyJz2FNxA9LXh6SrhkPzL7B/7PK
h96HMAcusoqtI2HGDW8ff/gScLihqrGS/7TCaEZgxHDP1ohybzHVejHmauJrxQqQRicKIJJQ3SHQ
4rSLOnsDglHssEpiZDfN9goiNFyigiQnSA91LeriHgaJYWvcUb4jh/Ign3asz13LyyzmluL1R7oP
2RqkEb0Ttjd9fdw4sMtJ9yQsNrGRoL84z+Pf7IFfpXN+zCSMQSeLrv543sRJHAXLnwnHEVbSRqUf
0mNmy7QiJM1tmkDoSSdPObe/heTb5MrN1V+QvQd8pkFE6lgSabZ0LlirRLzPvATaOJZKfAx/PUHB
zQhinRzJDcYodGUVtMvPwCtUhh4/QiG8C1hOKT54w8UNjDMI8comLe9rLy4tO24yl+ZphVv03FXN
kesZsmUlgS1fs0i9kafpPd33VGLG/tT0/0aRTgkxs5m8sKx7ARq4oBwWiy+c3nNADUSM+852npLo
t7aOQcNkBKx7eefv2Re+sJOG8dLni2dPxKzxPj677U9VRdAQYL3RdG2mX/s++F9AHXFdiw3+rnW0
xbR8Jg+FqCKT0QPIZhV+q+QclFBhRjAkvTCqHdXYVTsl0nlAkH5/9anrcmrHTPxGsjR9Roe+MmEf
GVk26plgVOkSa6ZzmL/rXPYE0f2YxE+DyfVqjVVbysj182RFIfBar0VxEWpyCJ1n10af7zd7jGpM
LsG1j6NOP6DEtqpC7dqzpuec6+i/zk3Y3oJcRXezxjwFmFkbgMVIGhey6cJOZpRTG6ENBzz9GqFZ
WDsfPsgS04PWTRvDgLg8ZXnf4sbQNC+I4HqpAN8LaR8BLuTwkhNb3LusjYDd3/Ohs1kMklRHOYf7
cWMzSAdEw6E1xIn9dL99aNS6CH2MurbX0Turxn/TF7ipDCJnUKIzM59eeoIH4tQ+v3S1eiXV7XoR
xx9yLfBnMEPxQLXviaTSmSjsj+hEi6o5/TslddI9ujHEMbg7hJfxQojRm7aZ1yS5dn3a/zYWiQN9
n7ndjz2V3lgw2pi7ZBtVK3sztjnWZQu6PTr4vaDYqWTpjMazYMtO4Zo8evOHayeENgxR6jg5t66w
pdCLme7wi+HWMuUM3jzXWE1+3U1UnM1dTcBg9miU8eclccflz/puAWt9xAIeWFBUaPTjJaH+oD/W
uqJ5PymBJxgxKpBX5wdZohCHtc+xDXayR+sjP8+ez5mu9+en/VfiU1h+ipZO8InRNcZ18hy0EqM0
Vg9XwhuG66btbwE6ZMj9vpFIOA7iXUyQhEp6BjEJNxoV/V+Fy8ipyu7qfg0I5rVv9dbCzWXZ4luP
XvCXM5HdF+7kRdiazjOVSfkiadEZrwlCInjCSltP30CWBHEd698vxjrYUU81w8G/9KsscHEDO+1b
LZ85JbRabYlP2nplQe+rTn2Lnc520B7/csuyTWtyKtTCK23eUmtOyqezJAwpY+Ct0Q0zTsuwXH3n
EnQhHjiQxr8q7zgMU/7pDmTP4N3vBOBOBcfLhNj4TV3OV1AEi97eBZXds7331IimEBYNNP97QXlS
y6Q6ohDcFzUouF91XMglf4hexUvgg+oLZMKjB83hRvtvzLA5/+C76bcBWZ7x4iaQjToZ2z947QAk
pLsl5NyIf6WA06BcMP827EJ//GanTGaiYmDnhPivYgLYefiDARAHLL5i1MjMMDLvscU1WRRPq7/X
bpT1tkI7xdarLIpAbxGZHf84SasTW0pOyoDfXFLzrOTdQJgjJFAVPS+lDp/AHEW2Anpepr+GT1EO
7DC8MOtF17r4Z91KBy9mzDcxHLjJk7bU7lsuBnRhU359krgLSlkMH1A1aJaNOAWCXElRdOXMuPmT
WrXrEK9DJ0FN/VQeIEjb6StdQG/3KRpEGhJzNwETuQS07thj7ThEHNjhy/wDRTc4QuXMGL5Az+Ik
BEQmIpjIInNyCfbiFeS+IYRoWascr4Dq872xrywmFoRWPtxryuSUyNyDIdPOEMwtqBg9mh7CBrsh
TgSeWHf+QDkWHwOf6/NpcZqgmd8ajOW5n0NJTWfvouiIw/zeFkzFtz86wBkICAgkWPq+5I3h1c6w
sP7JlAp2lKCxBhwJ56PV3sjiMPIGT5tMB9PZNzR3YGfpg/RPpdoMGQxnlqxiRwiyeAd+mFoy3CUJ
ylLUgdY8t+it/+PofVqcF6EPD0UWcxhIMIuS25uJCcM/ZN3EOC8h8PoUzbs+v3xx8e4ku5jAmip9
qfwKiHFhOn05t57PrzpIFZe7rzWM+KrdZlF8caoN728MMzoqIsykg0i6OTW/hax0UgX7cCzPrxUF
NDBYG+57ehfEpldQIbwtGdJ/qXAPMoXh9yHuy+pN1oRMDhf6oWU3B15SYJF2HNXOojybP1I4ISF0
1Nepg4Jk6B3POMNMaNeloBRN5OIJUTYGv90Sz70U1OewnoGB2+wVUsnbROS+IFfdze2XytvIi8Dn
BB4UCyGS+UmEBEr9OeltiyS5lLUwcr4oQG4CExlO8vSJ3M1HlDnXon8lt9J2rMWuRoEu335DAZcf
3+iKU8RbvybVUqWLBnQU870y3gIaMD6Qjtfw3dS04/vtVPqTU50jyRwzdXgm08NE6kPR8cRGFLiT
dobziBPpIGdkYv8Toj1Q8XOKgERyn9BeT+IwWVfhWD6jbUcb/220BMw4hW+i9zOL3/U3KUSzxZvX
pH2Yd2NPDxfrjODF3Jw8CdsaFF/sVaRTd8xudPEKQfTuwAA5hoYUqcUGWPsNU82zO97r8/6/VkLq
5sqbYazsOcWnZjCajLe3Wnzlxw/BLQR2eq3uVftkfFbTGtlCMgzPno29wgpTS5ND56DTBJ3RAOC3
r3zptyaPWfvn1MIOfW+4j+hqtzQgZPlaqwA25aXbftLthXkcCfS/9d7hp6RnaFyAVa341/d4LNII
MNByfbrnEcuEiR48r4XGourEi39pyFni0+4AE7o8YiDkYpo5b/mhqpSFbtsz4VPgCeWkdfLJwd8x
KsbYPo6iDdzdvLUDG4+lkYfBy8dBdT2VDxF1dVLQKzO0u1g2I9YsWylqUiAUhKbxo5hHy1TnOqKM
NHuRGPH0VnTD0jVvaJmmrMQjJxMhJ9GovoIKU+I8Tt9edacJfpwK7mapbnD8GRYyoMSHrw+gW8ig
atx3zhxfzd5nJJlJ62m53RjW0I8yEGCgfoN56AOhlYfNOQdKRk4ayYE/5wWBCEiwGvomeom3E3SQ
lWcy5/A7YpVsTxyvAscT6uDEubhmwY7mGsi56hCls4OwG0gkhApxVISqz8d9GgXTtQAhQQGBgiU+
qOXt37mbNAXU5sH9r7jH7Pa5ypVArNYw3GLcIFMFosXFDk0zQRqjDFmJmqFOENef3QlAjQvUHlIS
KtEz6o3zxNPJWM+xg1V9NY+DK4570FR1lHHDPSK1WZ6W+fv3GZ2td7udD68H5i2Iqjv385KpaV5h
yfZ3Xd6u+BWKP44B9W8Op4CpTAeFVpmeup5QsKvreLy3pBBEUDHYPCr1VgJyPRmOhIK8nRkbbCrg
YWvPeArKjhcfaZZ6CAnYgz3nGKSDu7wiUvsTWdlu0AU2XRzGe98R9XmNxOl1MwBFmwrORUiIkibM
/LaTo/tSEO2dz0PIUhJFtKccbU+1gvu7DVFvepznFf7b3d4RfhmMAcFNxtG1Y6a4lwYJc7tbMPWC
wpS+Mu0s1+t7HfJjp5Trf1sotDgF/aLkJ68zwfIquWfTcU20ryTb2i67dWpef5kSRQwpfn3QyTnl
Bex+AF8hu3kw6WTTjRcqrp6XWfiiiILWhQB1V/nSsMliXUMqwZjTx2JPLo6Mgxq/gSpgeiwRCLpE
RvG99anmgF06WiIR1hW6Q1eoo1kCFADBb6FsoSDTM5g86kZl3hC7syKqlN47Lm9/LAF3g5V7S2VH
4aVf8YPA08uBECPK+9LGE8WQtVtgUq0nswLcRk73x2sNMDww6wzWDJmpfNIt4iBVLCq5FYU5B9Xf
6FBYV6jsBii5iR3bhTnOqyapzMr7LhlPH19k+7/RYgQ6+9FPJRKBcaRxRmoSgMOiWeXERa7VcMkc
kIpIGn3p3lW9ljE5BR6cyh+RfTSk15Nvj/Zy9Z//8XU3PwvLqzFJ+9oeBQvTf4ydTv0ob54I1KLZ
WGr8TlNOsLgyTE/HN97SaHAUOCagNIuX8qITbSbs7zXpT9AL2ny0E6QWKGKTZOHO12D52ZtSsbX1
0IMWLi7aeufuDeUNgYXezCUM1qSRheOEnQhFgSd6D/gAIxoLiXzAqlXDGkM0yqJv6+zTWutJl3m9
kqC2u+O5i1Z4AETV/j6FXZrOM8DHEUvCua6Axlc8BLDt1KchxvGAv/elOtzkI6XGAPjYiGJPCAwi
hjeG9z3Mn6rUSuqVFR3ls/TnzmAnbcQU9fnMNDcJNL3Vi95gjeUpUcOTNDNJAFxbJ+tdttpVhISh
ezKI4slKRyc219BXnBAU7pjUHSa75OCbZ2+AwdhHhXeYN5gtIOdXHfJ+lboY5LlOZGH5Tff7KkSJ
w/VlzGISNucui6TUTmFBkaQRYkp0Dm3c2kB1WKntTMBrqhW8JqGjDij6K6W8Zqu8elTm9FbCbBon
SgU3OOCXsfN6yE8OJBNYHgJPCMd+YqLXLgwR4FVf83E1xfNY3FgGiIDIva85ZV76Kee/AT2Ty8J6
9PNTlgorvH+ymP7RnEeqPRvShY6FVWstNVteaPVjf99kOZPE2oMeWxXzOz3HYYfblQYFt5NPfD3X
kju0A8i22mivwDfaZOhc+J9db/tAh+DyeydXmOgNnVfijB3N315+jiJ99VKRQ+0y8vez5bqwPYo3
vF196BHs1iaYYwM3WoTcRhBIihxgvsirZWLxD9I89mh6leB1smAIeipbniLIgLY8XAOMn66nbjNp
R9qtnp9HSoJrqZdA7cDgF0jIVPQy0bfPabGtkR8GYEE5GmwQG3ngG+xehEA3pHmA9+POWIy6NZrE
Xgz2z0tG1en+1k4WaQ2CUswu43320xYXlS1G9YMyYf5WqOuPOzjGrBg5P/IUZoBAuWPsLxeRv3+3
C+a+1tMzhumRYndkVf1qcI6ntYTD0DBcGet1FRXIzFX7Yx/XrLqViIs7BSgasQAnUOkcHyDQqrNz
Vo+xbFYLTCRdpDKr3FVAWmLpdmkiCdFQAxolXyaqf+NAjJgd3Bmw/Sc4KwU5QZ/tOGQq4VR0EZq9
cfO7qImqGLJDfJoriYtcrAUC2cQ8Uuw8FNBRWXECgm0Welv6Xly3zVJLIcWwnmEFbwPxwlFz0fa2
cJgoexsFprXxHDGS5gji0SnW9GnFWKvCkrtO4KQ/RtlOFrr/lrY4+gkLPL9LfiZoU+a8dIsIyCAY
hn+RAzOoK6+zGlxcKehF383QVzsizGLa4DjQ5vvn8EvZ2mpgryX5WLhBtEWMry5QFHnOyuFFnL9l
DbR4rkt57yxNsImmWsF2Ju+Pybe5HliH9Sl5Mns/z+FUFof728HOZvlNBe749VfdMXsHmCMGxJCQ
oNsQLh+3FJzb51dQIM6vPL7rhFzcRhc0W1L0DmbmZS25lrkD3Fr6it7K8Y+dfRMutLWHCL9r7uXT
iOIAO408t0aGRjVq/rA8I2Tni1tCtTgMw1YW61cRnUP2EdgXgtOTNMk28WVa5HL0I3wHraLt8w7I
bXTN2a6bnOT4d8K8f0tAKeTfDTd94AnbzpJxJXfkaLefDS8fA11fvp0Sm6ypxVvS/0V/5/z/RdcL
xh++q8vCfw0VpcMFf4GV3wVfE5gHjeasN+oOtH/mleDCN6i0S+J4a7Jw4jfjNbTIuZfDTKqTlwCg
j2I5kQO0dQi56EOeSv40xcYqlJ6WWuDHsvR0H/0KLt4uq96XGzjdAXWaswukySYpdFSAIf69BbcS
567jYywVP4PLoVaXUKU9Tw5fwHH2KECXh0KcKx0T/Xltzp/hyHRxstxd2AOadUqEwfbSqCKyZl33
q8sI+S5B/qV760FVzYxy8yFauECbKBhayApzHqCOABA4Z6uqFhs6CZE6JVqk+dJaJQs0P19BBkSv
RF5ZVTtCA8p69X+MMYdun/2AxyYsZk1kl4iVRa2yzN9CIIjhcmHUzWqXOEbSKkw4LqmUGUnLeAdO
GVdINk9B7fKke4F0PqMAMCEk4VI90IMMgCRDHrXNu9gpHbOmhTAJS0co5ivsY6VXgNZbLWGNh2kh
VKfJiLfIoMWLKKxcj76E4gGxWMF35wnOzqxEwXC3kTo472mJprPrJZVR2UxCfRwg/BCvoLtK4qeq
Q5/cnO7dNo2cwWfw8IVp8Y9BkQ4wVC2D4h8fZx1RmCunVuxzRXXCtkM3VHXt88+WFNBxOmsqaGFp
CMi+VO174AVlpS4AiAIsLQ5MTomQNu2aG32edAOHzshEGI389i3njro4Ycb0J+c2F5nL/MEm+oX3
ED93uHt7Kdr2IKKD3fJSx3BJ1wHvTKto4JyQR3Hcpe/KWK696zb/cr66/6sVbnmpeT3yD/AV5K71
zsaZLpKNTcr7yGCNkgNc565Bm+NnBHrVNzwrw0lrgJEbsM/aZXrDvT1xf1HF9EchltxhdVdSGqTl
1jkm/1WgJHzCMLFwcS1UHvdvh/UPuwZ1sDjxkSuTmGxW3S96sra1SeqyYAvv68z3luoZzA3FMOsO
AqK5bfIF6qxSYvWW/rcj4fEZN5vrdPkSNhP0S3P6zxquemHrQDqpHpfs4WZ+saAz+ZcDSoWUX9Yl
85ogKFJKS1v1rbd3G6FHcD70/XkILCnmIhhD1/GjnYBmvZh1y8MMg/7s2fnUbAHNKayFvX02yy6t
kgYPpmXak6Cnz7t5pV97w3brW5f2n6XTCMWeVkPYqPIzJn6sxDSXYdeNyLHYHXEa/2H9xY6hAkY9
ThE9GcLaPivconbaMASr9RLEB9YRjFU27Pmzu+dwTfbgGx/FG9ku3U0KXDjTPg/ICWZCv1iNmv10
LqNf7q2lbSmc7TyBemq/hOdbB/m/r0jgV1lVG8KJovAYwskwCTfCccW3O3WDEyXrgRZu6ohOMTS7
ga4YmsNJoknJQ1QE1KAsyHMHenyxRl2PFDtFwuB5OJEI1Uw77On9C89mlFmVmuWSMKdTrzHi9/pB
P7D5Ht0PJkcPZIFaVNeBAa14pi+bNiIMjNkZ+zDPS1yN6OU1/zCl7gPfQqO8EdajQ/e7RtUvlRYV
0q3lAbfcVhE9WSe/7i4jzP4XNuG9IZvkkQE/kX6MZzAe3j4EDa8W3weG50Eh/FBNoIX17/Ejp27O
x0KPYNJXcQA1KIoT/p8jREZjb7i0qnx1pS8TcM4C4YDhnI0PxUGfEWAq6TxVsSitm52fYwGWQ3GM
V3OVzPqBFShLdPeYcE+Cf6tmHbz5n9q/XTrWVO9LHv7inuGMGPEvWlc9EUAVlRR+CQhZKnIgZMxg
tqFyx78+/5ajchvbMql5UYYV1FHbCfhBEnVBFcjUUdN8u+vj9wgXqGcsEdw6UNW8ZJ6RqPfI0JER
Pns/YpEcArZsm5LI5i85EcXgzw3HE54QrUUv3ceYpMYjeM4hHmjA9C/DiH22z27qlyGxZ1KTv/aG
LWBMUG7bcBPr9UIBXyb0L4Ean2KeJ2A1bUkekyCA5t5au8LIam1Bs5SARQr3+k3SeK8le3FVDmhF
nENz+bDecsQcO0iL4jJFLnOQMlxGQIYbsqTyrzwvJ04ESIEwl6qLvrwdnsnj++N+TcrcisNApixG
Nhz9lfUoBIEwiDt/mUrB+ZO1Hp8khOO0nfEZCW1c1jWBGmTM8Aoh4wn3FUzfY0sv4Bvfev6nriUP
3+7gedg/aEl6Yt23inJLLB8I81Fy6ZFxHK5ypIrA4r41BDW2u/bKmBEL1ntwIiXGeoSNoyW3O5Ks
YmnwBDL9oHj05Yuli6WvJGQmF8mhsJJ3+yGcv43NMvZtT9IzzZ+pCDdLnHfAYztgnYWvPISB1acb
DM/pUwMf3SEmsYT5PO6WwICW6JVjCZHzwwUhavbal7L9rPR84TctNN2n9lC0jt2orW6zSwTO1tId
0wX1z6Y+ZTZMFtlNe4ZH2/H8AuXZI4SD1qUoOK2EwVteG+qBCjZXyObUzJbPypvw8yFmfHV96qgK
ASDEYCsWVtXJ3BW6lDSWM5TLW+qGD+qGYamVdRQu5C2vFD8Esn47dCVpOB/ZkUyEaMqlwmorECX5
MNqSfykOvRMOijOcJrqGPC8VCY1bbUfDwdCXGOr3f2GwWAwgp4YyTXGwRtP+W94jzxjdFMJupZuI
e0JjO0lukbOZ+7A/uXpVAfKGKdihxOVVW95j5PtXjTL3BCalPe74dac7Ders6TWCHp/P8Kja51I/
+EwryWsM7BhUYyigiF3aFoz7vcV9ETz3l5zyEVoky3iwDPiPgFDWI72w9/nFAGB9GV0S2XhVatLE
WVJA9hNRd5gHIRVxeKqgmhros9tFbj3NtcGLpmmqJ8KQ9fG7q/6bA9+VFEyGLcr0jIx7g3Oy8tmE
Xvs/5GetqfHpL16MTWoUcsnQsyfEk3qNjQyuXiMRcZ5TXW6CmCCXJYe9YM3VYmP+ohoXSRvL51lQ
cDA7y/FBmprfivk5+i4WShKXfdxlwPYlh2Uq5AVD/EMwnl4DX0ylvEP0GW+0SEz/MW6jMiH4//NM
oZC/WRdVOVQ+KZ+UXntdtENnkvgodLvFix5FQtesK1bS45WfNNEc85uzyu5UN4hNQ+YiTsW3xn2P
x71tsQ9/1L1Wy2L4fjO3/vfrcbLBC158Yg6jt+i4jsmiA85zuydCBbJ68v7MYXtdkUzD/ZCqlgg7
eWySYzcsr+paxdQME9soiVES/I09B1sbAIRLhHgsyCiN274vqW0ITHcDDMizTizk4oIaOgPOkf4C
lW4xaBxUHmzctfa81qtmGHY5Rl/TQhaUIdL91vgWe3prUs0e9mVQr/MWjT6ChCJiH2cCxiwJSzWe
MpGBPapOhSCASjd/Y3p8pFvOA3sKGCtgeiaw0KM2+rXv5UWgk7IA+ZaEIET19+L9B06oE001NiE2
gUt6h05lhkOoWIloAU3E8SLPg04Psz2VVtDQ2Yzl7luGBZULnEhAAcTrFN1f9Mf0tzuceJqdS5IH
qgJoUnZXTW7RTSWooj1mug8Hnm7N+31waHizJtpwayrbpifAyJWQC0Rt1DOgYDqBqoH5VlqW0YZO
Wqz+GMSwFSSVWSlCEy1F1cwiBaeiqUq7Z8s4mzvq/lfIt2Yk1PCCdH/jLdOpbrELKOppfkPNZLDN
qH2k9qHw/OZE4nKQChH5tQdqxj9lpIlXrqZ99waaieYkC+5TUIWr41gupkqy3izGrugRRYPpKSdz
SDz4lnAbSxdKFigY3lFCnCg7/or5cgYOVk/ZUnCRpFF5xsBiBVb1BwamVVGJ9ogrDk9rswRs6WdI
rVTxom7gKVbQNEa62vsGdT1anaQUTaQVtXBaIBt/YORHm5juDcCyRlPILT9+KRHE6r42TcHgHQW8
U2JVafCXzUK1O3n/KodiAfbiXnY3D6YhjFg01XNlmfpelSwpIPK8+wECdJ9a27zJKi+Y8I6rbQLt
x2VO7mYFQpHuQBoNuVZ3A/3egmZc7v/kIa+KOIbzoFrh+ruAjkbldr+/D93tdU0p4IymLCO1/FQo
xGJY1QQzPieR8nzgiYLdfVzUGw6NUGQAxeuAHrZuheOb6v9x772JkC6sgOp9B65BZ+VrdU+XajIf
0KoNiILztGBSMecCPmjLMTzaKeHRRV2PRRkJX30w1FBSn4stwrqKLVpx/7SmJfHMBh8riOmHipNb
QGmIYY1kkvphfrfXxQRGv2otb4USqtJpgrVLwD8+2DXnhJduQ9uF7goTjKWOfp23G0nWD3zypNv9
OpyQpYxKVAbW9FbybjlrrYbJBmbZEfUAbBP8dHEjoEjlemBD0I6KkQeuszkmB2xHrnMkgT1uqi9g
5KgRuImu9QOvhq8GFI1EYHQB29tF62mU+dCTb2deX5cN7qd3qQFYSP4+D3Zo59qSOCt98swVlgmn
9H3ByVX48AX3lTB3S8eDWqktgnGJunvKzaCDZGR5u5CE0MbDJ6VKheGW/ie/PoX/H7veYwqnsw7u
XVaPx1/uP1oXmlY1IHoen+F5oqdhiLheLaekHp36ckMQ+1VFc0jpXetRMoDERYJKBF9m+mSyfSqR
Bue4pWpNhE/wAMgcJagLdpb7wMm+qouSW8B1VB6xYhZXxmGQxX0xFcEOPSzbGIOP1N47ginwrwlI
QjlQA7p0EOYeqcwk6PyRFCTtxoXPlLWLC1VDtqKmix4LkYY8sOdYZpBPDWrx2ts7pJVb/LRflkxR
bxRe7x71cVfhVR3ubb+Lc5wzzMdOacq15oMCptMFQqNtP7/u1XMbiim7LR8pauPaD80ZLVL48J2x
mmtLdM0b5vKmSVUlUh6I6kbwo03faYgZujJooCol8vVDjtWQXn724ffBoL2ls/DTeQT7j3Uiu5N+
ONS0qMq1r7bf1drhDbm9LSh+kNcJHi1dj6Eqw1iU9x2A9oovliG2+hVzjlcP3K41INhfR3BoUsCW
pT9sLkuXvMz5MHvjCZ9SBnrE2Q0VTcQirlYJQp0bJOhbv6gSjIml0J4ZS5YP8E6AJQJfbXkpno7M
AkwmQ8UoWL5utLlxlYNMMaQ9cKRYFfboHClk6X3mCRGPPgiddz0GgXXITqfdxYCjsFos2Bi6NLj8
K3V+DbWRQ4HqDrhxRX4VaTsJTIaRmHI5p1kElSKVTDoUsOajW/Ndv+ZBhv+2S9tvek5ZLShhfjgs
Pq1N+9LFJkuFhYtomJ92eyLG4fnw7kzohoa5Na5ziV6bynptkQL5uc3IvIBbyrUlsyKILFkUS2X7
b3EQYTAcWFTN/rQ8XPcFjphmTHWP2H/cmaZvva19C8afGL1O5qSGluZxkuxAQQzSbYZ8gGACAOp+
4JsBmeF1nB8SpFylp1NEKoiPyyHkZOdmQPHXQONI4SgDIsoQmDemlynPOdBoDhC3syMb6/JypnAi
9N851aVxJ3JyVBnZyOuS+A2PmJIsbu+rgBPDi1AQiG/b38irx76uB3MaCz44BNK22vpmL9s6ATt8
NwB73r8aXHTynkK9r0T2Mp/AiAv1R9T9PwTPIRhu1dcK1XePMdj7XqPC7MbBSc4XNKmXnrH/KA60
1Ts3SBmRqxslfz2tZAuYE567mxO567wuKVdR8WoapOWEHw54X9sgcR2LGIgYJ1LVMAUDRPPmcWvL
z8yaKDEg6iuALw2xOgTsAduzwmMu1xonf+vKP7XG0GfG/pCWmheLOYgz3It5611Iw4B4lQBxGAJ2
iqPAkjP5rbTi617H/f/6XgFUkvOm/BR9wHU9KNmbn+YIOVoL27wuqyl7fMOTlaKNkmUlDs7n8/Z4
kbeC2WuYPCWN4+Gm2+hsKgLmAChSReIqAd1nJ4CDW+Gl/FUCqUqYZ6CX2bvOCSuCLUA6ywDMsLVR
UK7fE61AFx+48cPnclsTYib2PTPXjrswoCAKCwsbOKqtI8Mo3NgTCoTH8WjxQzOLvVK9L5PLJFod
vGSNa5vXoT+L41dHVxvEHcLBPwH7NW/RgzEYIqK5SUmkq//HGQO3Y+M9y43F5cMlTpDEJlG/zP29
klc3XYnLTEEuXfs5zGcoPqZPynQ32SW0Bn5pCymB6R67ZKSHZDaaZ4X/ikZkQAsbOPjcfXRq6TJt
/hfmQM6wv0D4VaQCre6CSDNDaHynMitoHQTDxZ8ZslvaXcJ2Rr2e0eTz331fXEXiN+fnF6J7EvG5
FofeD44tZacRByXcTJvaVaNiPFUA/tjipe7JroO3x60rLdT8kpbRa7MHmBFkctnJycR7e0S6w6um
sMjnY4McuWZY3fE2QEvsZusXl1sfU+edqm72S93dHN1D+UKLUrYziq1KlkHwRbRNOD14+z7ZiVQc
jTwC1GaSRBjaU/Gm7Z7UHtB7roxROHSOT+zHQ2F+U8K/c/KquettRCUr0Xi69seSfuY7tcnT+/jk
NVyEy7aIu/Gh+effATF5L2g8aKvXSp55YgRHxW7a7GVfYHBHV8h2tLgo5DjiWOg5VVz+sYoF2OwN
gst+YiYb9EtT3nWUj095Gfok1mo7TALzZvy9j8G4HWgvFrFnFXUT067PtVdVBpNMAyOkoNK0gA8M
ViL4rmbAbwqmfDovJkZwKF0i9ZF2h0kMxazbP59YFS2CjsFr1R+8nPmiVlZx4SYTuZBgC6X2tFC3
txjarrgMzEytG3L3qN5yrgikgOnYiS07aZH4WkqyyAuxpIapbakM9BxWEvsq7VgTyC0tTYc59PTa
nf+YpoLTUaXM+KIEnjIzqjIvJ6CpyGe8WGBUpFJk43va5rYuk0lzQBcnGpmnVoCMWAKgthVgW9+3
nh9dNz31JUtX2MRRap9fvw440gjPCVHD6p0u86QhoJT6+fHrQVatvlzR9qXMPJex8+k/w12gSi/A
HmBsP3Hrj3YsZdp5KZsuxqKC5y+5vEgRkYAWhHyy5TDiIOB+U/PRPM6K1kch5E2v7tazMgWii5Ot
HM9J36pQPdVaCAZOLONbvYcUAJdag6ZA+AgvAY43MF5VHhnP5ooeTyBTmnzFmvnhJBm/k5Yyfrba
sP4iLe9xrxE2pwMpXi51eIqUgimmShyfUFqYvBE+b3Few/HUkH0XyQ5e4BGgMpOLv9DWQynqCVeT
T6laqERwjFuJqnPvYTNi8bbb3jHOOM1m4GQdrvWEu30HNUsnmKwxc4hlT9kdgVWaJ/4mPOpWJKpj
xk9HKclqMAF+DAdnI9y2IBtIWEhMBRWnXYQvNrfdZvZDc26p1kPj1ObLoVsemDl33sdmyOXWmWAH
WyM/+bSYqg08Mg29+IWbP49FomkMBikcnZyKJWb4HQ2XvvQ8hLoR/PnEUZFMjitGi93LZjK+Ng1j
DlMv5d/VhbWCptFsPVLk9r+rYzEXAigG1Kf93UIzvNfTR32hSvHzsVZ5wsYU5theBL3L3jLIcGFk
NFP0e0MBEd3SBYCK7B32o7E8jEXp/0WbeO1J9uruzxwoTtlzSrJ2Re05FaicojPIKrf07lFqaDSL
8CXgZuQAAcJV4AeRf1nExsINrbcKeH0oxi/jAv5IVC23BMGzHqRiyFh3VFwWAaOz7LfTDZttJ04V
w3ssFDrxQnhSCo2c1kCMMKpvDIustZaSMDJ6Qv5YNuw5vP9RCBAcDz5gKXGHDjmW8ZM+HeS54mZ9
2e3xXlUYSs1VO6eB5Mo/RXCRYVzB5yb6pv/k2Lr+gUWL3fC+PpWhtkNEd/qoGqFKeA69BQJNRh+q
PlZ41zq+VAkKbx9gkvHoPcbLrY+Mp4GM0jPY7JH01+phpiWCx1ziutt9Srm4GqeGFTrb8Ryoxnu0
94zVqpOPHJLki2kzNQlo3SNlaWN//SjTwjrQn9YxxBdMADq7mPc19XGRvMBe372rMYdIYVPcJ4xi
bmYpKTT1TG+5huroBkHtVPzi7scaxwMBGxe4Bedd66ptHk59HTYZuJStVl8BJeWcGRk/rNJkNT+6
fuTu3WxB0llmcBgmvkhz4hYorbPEtk/HF4fRMkz5nNNX47SeRyfktqGaWarw36vu/MZFA+0Jpn0z
Gj19+3VMvB+NzC7/AcZc39hE76grGicwlRr2Hr1exScoUO5TeEks5Bc16i8Ni0YslpYmynN569mE
njMXXJySom0jM6aExUE0DV+IXKd1J8w9UrqMZJU9RDJRsBg5HH8zftB5zvlE7fWvRPRr24Y84RPR
R+GGR4gH5XvXtZeMlvbfIyp8CKvziL5njh1VYkH4tfPBs6sMbbiDwTG40C4iGyQrhKpsCfUtd+W1
OeAvIw8QN4zt/yqOsZ4SBoO9rCj39G4GfMcXJK069iLNkYos+emAzjaqwks3eOMWifyF6oUvDM/C
kkjSlOZDnhkHoe3X8GMHvGuxP1gctJ31UKLa26O1XbqOaSyDFUiVaFkYjeHI4/GIwxSz0LbFs8Xd
IoikJRJSSBdqtOzKrJBG77W3P8ieayv3pAXZnxEZN/QSjH53T5nTjq+UN6AHpZislkN3l0FuJtTW
Va1OfsV5p4e25F4bNJ90ogqcm+prPyigxINwCZXw8bt7ymydPhjqD/+N/Evlh+82xo8uwQJ2qefS
OB1U0Qx1EY1aq/oKnS+OW4lzW5CgdAsquRpar4+IwnQ8SgQ3x4L4srwlCqRDysSQXQ5R2EeUN/ML
PYt+L38tfuS6ClrRTCFlYuOZvAlUO05qvlEt4AZoFLOsUnAS2MLa7n2zjqcqfa2qL41BGFmOvUMi
F1e+57t4wKlDHYca3abD55WHa5QSaY1wIiDDvuu+GUcYLtGUSqyGqMTpMxLCgB+u+Hs5EVVFAdDL
WCghSJt6irGjBaOT+z+I/bBmOyBt4i7/pkBFSbKSsK8LDm00y/NiXuRpZLqd86EBrnijhVSE/vzw
96127ockVWZk5lZtpeSV8ylhYEV8qOifxprqvXeFMKmMDwRPUZwwBlBju3lISveFPkgiaWt3R1RU
Y+ufS+e/RsJhuklh7bYKc109RKIRWnQUaEXHQvYxDrFiIMwpQ0p/0uuZjikZ74kkFBM2EoF0h4+X
nMiPR8zA7qhnvY9F+e7D4wL8/idPPGYi/DfaCrgoGiU5K1n9emUn9IYg8fcvM4ycpw7ZFKkZqkY8
RrSJUtvT2n4sUnsyej2wLS/aHCS/84y/6jcAy4qDH7pE/CXv0szDqakquOnmAbfRoQCYGRPEgswF
cGMhVDDqPxrPJ4dpTTNA1mC/Q8VzfotXe15b0TOcm9gnUy5sJBm7CVZmERdrBBLCYsN43mSoFoYS
/B5y+0Zkm6ZtK8vbM61unptrC4Hvb13hf1+5LdNWoMsPT/CVNq4qjHJU17IMjvF//0qxj4BOnKgu
OUew8xS8djhpI2OXHq8OfORQn4VSez9UxO2XzL5mN5aHaJ11XexeK4HuUoz7gxa1Ycgu7WpmYnoZ
O4qOAFQ11+Sa+IL/NInJIKferW21PcGbCSZrkoMPzRZ4ltpsIsYTC1seF4K68BdgBlnZx5bCG6n+
eNR9EotKZdK1tXBWFwdVvJuYXUpIHefKDKUZ8JYrReZRsaPNmsXWURfiwLaqN/D7TJrvPc3TM93e
dQWAraMILkw01WBdHtp+x2lWyx3d0PJnl9wB9aS3geuDjyCLk0vlcEmzvcKHsfxpyLR5LIXiWzij
mNj/cXW4jUGfbzNJXMy5Ml7VrH64eMkTTQlY5kdBSuFK5i9odN4R/HrZJ4cKGu34JD1PvXNAEOZR
3X85qPObBVewhrzrfHFlJIp6sn+yYqrqENcSWTmN5tngwWprjSBZ2FD0KPR8moi+3/wsYrXMAyJ5
AD488eDTDT8U6yxMKggpxXEcM3VIq8nwTf7R9j/Fu2kc3VfVae2NVWTHM7a/Tt+vosg1HScS6nA5
z8sc0bdTqAHtisZt5ZyK++k9W4qUGsECg8liCus5+7a05zUEpto5cn5Yl7s88tf1aXZUHGJvYUDR
k/R3TGh2uTNNECtIeav5McHGewIDSptmktpfq63v65ddNEAuIRnmMUB6v98wuH7cvVlVzEAOJyXl
Dl8g60CJszqP+diZg2xV+htLl7pZ2jv9qzL11srlvWv7s3dWugwnt7Uhh3oLnubQvTLFQYJLsxAj
ls22ucbW8Qw2+IQdaI9SIGj2XDFAVFrh0T3uVN8bUxTn3ZtRaR2KQXn5K7zYlsl+X+InPi2kvzPk
e7qkoVFmE4hZtwmCKodFqoLgUMTbnuROc/cZ/9diZMqP8uu25zUmXyeXpaqcs46ePJIFCNcc6Qgh
78ombqgaawWxG16CE3U9YQiKJ9/syPa5m/bpIeM6MSSesEzV0o0xVAUlREJJMKPVE1H4hoLepQ8i
1DwJoDyb2RIx91086gTttMuTZkJKS654BmL01ATrrIRz44ly1ihA7ujwBXSQtTCsmTc9+wB5mglM
KtybYCMIzlZ6J5shKW74M7JcjyDm/tSOPTnaFyT9+kF7qcQGPZVrQX6rwYJkF6kGgMGmnkcUAe5i
hgpORj0rT+xHvjCdgP/IGJ5sWwN9RTnWF6hCl43uXMyXpNoulOkUOxpbVaO72+oXQx0b9UgbSb+e
v4rRqM4zuNbBl60G2CZFwV1j0AvWCRzwtjg/I6fBUthhe6pemEUiJBwLKOforYzfRpkJhqWydcij
8Y9Lnu/2vapcgArMKSVnmcTBKH8hbfyROLFBO2fIHXrK0onuy9MNkGijGc4YsSq9lqm2f92XGEv6
uVEof/pNXl5KqaOw+zQRN7j19bS/vjgQZh/9fyAFz+IuWJfzif/xY/Mg8dR4wR/rLracwr/q9pDQ
xf6YzK96fgokWL4SwZyWal67MG3k8TmkrIYkNJOZbboz/rfetetAnh9oIgDN6AJFnyHHu0CdaTSF
XTxEIaluRZ50CYlp+bvZQfctVTi/RnogvUylMND8FkWU15mfLtvKMdQmi8PPh/8MHgb3FyNQ3abg
BpW/VvGRoZt8ENykN22q6EbM2FdzSF95ZUhYuCb15i/cNfB1s9p6ddDuGTruF96NNlpLdM4HUffk
LY7+PI3FMpWM2Gl06pH5Sij1B6MXh6YOuMqH1TcmxHg7phOafE0BqPLvFWJHZMtxcqValSyhIJhP
OL35bemdYNtbN2hvyEHHrV9ZV33FK7+izs8Lia+0S90qpNwJ9u8Dp1IJCsF+6PcVpb5Op2WTS/jH
PcWeaqQ3Xh0zhmiJpqAarIc8rcw+Bhs3JtwvpXfxWQ+b/kh7WmfnUKMCZaZEiVjPdFI7ZD2ZoLVb
INcxyl8Ly1PQJyJtlvcTopeyN8xFzHAtLOKOUN2RlUqlIxLSaWjAWG8NqqYt5MqG1z/GC/nsdv13
R9uOngqOxjM/Q3LRxd0Y3OwcMcDI/VcttK9EgohfTTV/SDWfA8Wace5sepxJgj90ClTKP7M7QnO9
YeVLUOdTtynEejDAn3ojOFRjEEL4BZY/g0xv9F51luXheh8k2wM+PfzsXCI65qQRNaDK1deccdB/
e58YWxJ+OdTW8vB7SliYxizSQmSwN21DTINl8YRPT4Ph+Xul5YXw2eO03LxU99qAys3gcQ6hPURD
PW2HT/iyIcxC/Ig+vCZ94lCxNXNu/0+HUcXhqI7ryIdP9pYs8B8l/cEyQVmm0TjOXg+Wihb9EmKc
P1qUcswoIDpsPY7KJO6Yfvw7WQMraQmh01Yc+YA1RyCH31Ei8ZYpGedFdnCKAXkQpvIFmlC+9G4Y
GsbCygAscMR7Okm6y9H91CPx2o+u8/gUIWaPLKXkIGpYKykSohafW0c9oa76eGtrVyU9GzwJME4a
X1RaCAc0EmHqdIpgKgHDTLs3UUbkYd0Bz6uXXhMvCJKZPOqFhHQtLcfdI3Ler4LkX7f5/2lMJq1W
zSGSXOHnmPTYmYk5u5tpm35qXL9gp2FHU2A/E6iq1OYBD5NcuyZMSlDamHbJ6SjT555/MvXRtc9Z
VCmI/3fsG2oSuEQpzVPNlZL5dSktKsAI/s1f4uehRawvBLY8Qv7hqAtzl7Cg3k4nGXUXqwc5rPKO
I0x/3qxUiptPTRiBJxf3E4Q6V62S1TZ6c3lIU52QNQ3W5VfBAq0tbT1gTDqRKvRNBS1Ez6es+XGc
zA3JDoGgjyKebk5F83Zh0uhB9Kq2t5TTRh8G5tsFocbSAxn0szlVfhH/DMmjmQ7TmwHPXc0uY218
zjmmJEyFVz9cN/G+bARo0AloY/Bj2aZrUxnOkJSY/nrGWAVN/czXACreiTMe8Y33YBnYLzFLYens
iMFO0D9+4Yzj4vbuMkHkyNzAJYF1duIUf0imNy/ODYd8pW/n6iC3maKx1/jQ2zZX69K9ckYUoQsF
hPqaJGrhR/GEJWpHumz5GG4FmlOQwTf4EA/Q7nhHKhcU85PVJc54z9EzOOGEmxYol27S0A4N+Gfn
ljNXun56B+RRSvebHewEWE7eUBphjS9lT9FvAigFPAH8FUAayq/5EUsQWtR9T7s6cHQRnZNXCOaz
mXyIKEXwGna2qxE2Rk9tFheJbhHZIn+FphpA5OnKP0yFKvIenpH0fGs8zAhfjqpNnoAHS07Z6EHY
LtRsQYTYNOXz6p0AAS11g2PzyUukpUw08/w++XtG8bCTwnwOixYfjnoDYNn92yX00y0j9KjGE6gc
Ad5FFuN4LxJSy/iYTlVAfon59eVQR8NKGt2r1IdxCX3bRmfDi0fpcVVyNnrzp5UExeOA95pA9LCo
uroBJPWxZYjtmdMXIFzOpraG6E+lTbZQsT7e/lPf1dM+yvWGUWKt97eMoHVpodkB6QEQI1u631I7
it2c/yFi3LMdxjh9NoRT8lwxM9vXWGBJ8pvb3nrLafaECclo1TMSHUtc/OK7tQ0HuhnFX7JHbHVd
uCOwfB4zovqqu/+gnA3f0RCjd4B4sPVTX8miHCd9bFFGBGLQZApLj8w3bP3zqjEuVpHNkTXO4ShO
PPugPF9R/Ids6YtKvuL/87O8LNX9svFcGMik2ceNsbcEB9oRXTeu7eFlTzyqHBSVjW+niMV2tb8c
vpWlKsPdVBZ7icVLdVXex/Vr9/SQs5jqWEMmf6k7VXL5+TyoLLZeY3KtWgnt/IchH72oBPs7pQGk
6GevDRveZT8C4RXerPaGz9dCmbZsWdYJn0VJ4OCkCPG2v8UDOCJmUblfDcYmS85Y2cr5cFYfeolh
yGBoJButKK7mSMlpeVdTfxim0Bae+L2pvhvSWkeSWiqQDBYYfvmGEodM0wcfpNtz/JVw7tgEVPen
udLuj0fZoR4GqYvZj7Y1TSiYQ6Ju11WfarudYZKYu8SP78uZ6Q1X3775sQ9WaVqRZdPUYqzbYNYv
bW6ep1yxwiVKi2GPnfVo1cjHNh9HcA8ZW8XW7YQECMa/CF2TbjvryDNjSUdx4hiS8GBie3se6Uzl
2EkQHiJNCmgslnw7OMx6f64Pj71d7tny4QoZtU9cE4MdxTb1YEek6mNfAiONOsPFnbph5SE7GcTR
/wLWaJLTQHwtowhdrlt184eLtxW2rJGI+Al+PF3PQPEzUNEa49zGnoqD1cqlgvlMhFp3RHVpnvfU
RHvlCW3VV150TNhlc614JV8XM3oLTkAenMqr+9k5YvccVIkQ1VtVEtKNf7ERRmKr3sQFffsMoFLy
HPaOILQolplghvRXwmbez2BC/hKVZj6EqTGssQTbms1sFrCJ+3zdA4ngAbH66sYU1kkhZxTyns0o
IxCj+q/KcEaiPusWu6kd2qVpY7WjieUJCLgUGukb25eWiqssQwaXaFcvQsl2JHwDMzH9iebR8sfe
qh5/dfqjxJA3QtvHukgFcEpKj+54j42nxQo75ICAGlLOPcGfW3Fjs+RegJh3S7YyBSXGdjkWdsMH
MzkUlHMSWg5HmOk3woduupzgokD3UqdDu7oOgzl8paN8wul0GDLO2NjatTrFXQX+F+MkkWU1my3I
ofJY28LvXMrOjmqTyKvhDkEfPBaG1kjkS7hfWR5ZHI+df6ji5J2dMe55YB9S9/MYptUJhX8iDmvD
0u5HWIS8Wg/7HysToxO7FAC2vbGiukFwhVx0lbTuCLz7pRvCA6l3gBRluBDtKPRXS7cM5taLSx4M
pbhfzEG/rq30V8IIHqrfOqym4PxIAqc71w6cFaD3roW3ytwlpSiEO3k2wOrHtcR88s7laBfPpyWm
6yr32aZ9pg6GDrcSAz3/XIrwnLGvWd7P/cxd5ezemNvwUZNNtxWRVYcWz34JiFoMqK/9ncImtfnt
MK3JuISEmRBCSvuNA3dxpwltMaXMKgfSz5x3lpIGp0UVz8juJtTqkQ6KST3gCsaYY9az0/37zCHY
YvbLN0irXW27T4C6QeWeUw05lBe2b1z/ilh2XAsxy+uirASG8o0frl9OV+Ds54WTdr9RkQgxbu8y
Q5pA739aORfserdBOgXx82zehOZewM6J0SIwfnyI0p0k8pDTAlMiJg4I7/YI/JSpOyP4+XfiUnbX
YIyarElh4FBfoRNsHR9b4I82f1sD7sX71HbQRYXFvx+6Zuco/TW0nacGQMG7WrwwPLoWYmKVv/Vk
Z09hz05TAs3LRJs0pka0UPSxMchN++abytwKk27Mgl32/Xr6w76XWHJLpyQzrYT2/slnBe8+sKFP
HRfTXOa/kW/bjO1CjSTS2Lx9NrIarOlIDJhjXHQErCWVQnP9OzBUM5OUvMgN8nZ9W0OotXkSxCTN
TVbDEzRBNb6hy6/4GLgXrAuTGacb5uxvJlnmqvY7oW3f1hO+BiCJ68CE/XcihcUFvSDZj1cqENmw
u27O3fa4cX9DwBA54TsVzWlcv1CpXHZLtGKv7acTjHU8Vg4c3EfrynqZ6TGC/0H+y6SB3KvC0obz
gU0TOfvQ3/qIvmhS5V29rcAM82bi4g6dHvJTpizBJ/v2cawonEJS/YkhDHQBhRgNp0oOcCG1uH+M
9bnPxXhK4P74Bmr465B5FVp/j9tsm9MlBlp6FyxdKYv8w8m6tEPL7/qXP8vpCvy7KW1KIJpMP2n5
v/CKGHVruTTqfCrlmRNVqvb9cB+2LraisEx0F7gsd1iqx2Cf/pB5WfRmH1Zyi60fTyUzRS+FakPe
VuLnARQL23BWcP3R6wOCLPPJKoY+NTebZsBR1YH1RQqbB/aTUafDmhdW96nGJa1NziTDsk8zN1CZ
i9hAN1XrwN0gBQZxbBfY2BWWMewhfRJK9e0OlggRp3qdIp9MH0rm8VtOQ+QBDwcHjcecs02UGYfC
I79loRX3kUp2ZKbZMq/5CdcrXChOWJ8wB4vz0aepAHl0cUG61WoS+Cc0fIAPQ7Co4RYYHhT9885P
66vP1F5bXYZz8tBdTDSFLgU5yqJ3mtTqqHtsUV1U3sYCBUAuHdtYA1k+4rnQxOR/f1CcCT9ki+HQ
5XJtbmyMBblWevo9tVLvVbbUCPWVLAUIIyZDQ/drz8z4uHUQwIvdjy75P1qtzOzgpQQi2eeSQCPU
BN+Apycr1dbejeRPvUNle+sCrMoLSnu/c/C6ZAm7E71I9rmApQxftKFvPKT5g6UM+KABgRA5uddT
sIHK2W+at/xbmi+nyYnrRClOIFZLZJE9vVHyaG9l0YeKI8NupK1FxwI+PUAap2tC/kwFdz+w89sd
4K7ePu5sir5C4k7/y4RgFqk/VAVL1DjKnwz1nlSFac3BDDP0tzubW2QY8My1Qh1HzAncgCblAZhe
eD9saReRNIY9KCgLMVAxpJ7tpkSwMwBW5TOGWYbb8B9aFgDHVPiEHxkffjt2ZYcBJf0U5ZIqeUh6
iJRV2sF6jUzmk6cHToi9jcchTPNotrlCNvwWbW4r85D7plaCyTC6gc2TlCtxk0EOYwR6yq177gEU
vtVpMGxaAZuc7/pib1canWEUtWvKJeB2w+sMR9Zh2hxueqY+XPafBCDAHCiQ3DqOatL4dqbXT4Hr
iIc4m6hXwm1pQoXmE8wia7XX6EsXqcxKgkBdodYb5BhurkpMoJLv2lV2I7khzeptcDqPsYo08BhM
hgZSsS/DR+3ZEYdGhcjGrdYbykyKYIyRuNNMl2S0O66SbBTufG8JYGDmdxNlOBPcaZOA22WOI29z
gA2h6Zbt2/XOrNj6eQWPn1klRiAjJcTyi74Zzt7NMEY+H+JqaIQwdEW3of61jWamS3x7iJdF9bh4
eGPbzX/VBeaKA0cGfy+VDTuYUiBfk1tQO03xdb6Ga4WDEsxmGo2lsKnV1rUunBAJexm56Oi6HHZ0
3mJvn+K85n7l1WTYHr2/YuJumFMDINYHfy0COiIBBWbTKO9B53YeLJGCNrh/XuIO/MFh4x9hTYuW
fzLpeFjBhPSOOTU+M5VzIVi4lks/BzKNHW48vu+ZDZYz5pULREX6w8eNUXFTLUYnXokJj73JMAZv
kh57YDoYJDeVnBJSuAraC2X/ha8PZmCnmtcMJHl1MV1v4CRXDiITEDFxc9D2q4jCYaR8G3qnxyWO
dIfLq84XmehcR8Ojl81cqKzYuwRln36kuJpOzuoSap9mAgN/qbedVnT3svCQWBMQi+h6kMgXWEMM
X5F4k2+BreeLAOTHzYLCsNq2nxiiapBHbtrGfLdCjV/UNXfd1bopZcriWQx60wuPeFfmVDKKym/d
y1ZFzpmU8u+mBkdtDRDxgfsX8JMQRkvH8UDgAXN+oHZtlU/cM/cotHWF5gYo5MIe9ZbgAll4B0q8
WyGz7u50n5npHJT0v/l5xHTvIvcuePgOIbE/Vgsagj+U/PN37x+E/sGFHwxHY9p1W9hYbkum2xlz
FNLbWWSL5RUiy2BnjTM8B/Rr1XimKBw2WzUpO1Sg69oZkuESaAq/QF4t01NlTk5W/Ba/0DLIchxS
dKhUfQRspw72pOy0OLEisLfHTtmLVWE9AKim0k59KnJNJMgiN0bpAX46xz0YN9cDss9yYPWlxI9s
xmQPE4RTaJVjNZyJn2PpI9IyLq5aIwwAVNzro+egPI4Mee4eX9rhaczYrqHbbXVTgHm3mBPTmqt4
G3Y1zvo21HrgcO+ZnyGRIUFhy+Ww6kOpWVL7xun87IX7UWysYaOY1+oos85tnJAQdrsP1U5gLczV
GaI6MLtu21obB8icSV6XSe1BJRlpHSuC2aiIWmjBOilq29VjaHrTldpTAY8OORyxcHcZWiUINdWp
bNC9rOctHuoSZjM59zoFHp/GbDa4Atqf2GI6yQf11tax8SQACNrlcJNcbqsOVNEbzHz5Aihi7ZN9
2UBMwJ0SnFxbwIjERKkFCs84FNv8007DnrnktnnNW+lYrSbrMWeYNaGQ0NCSPmajkSPV38QjlB45
acXbtSFpmPA/xxghgecOUXJU7cgrfTubnbF55s/pbpGME8vcjyfU17SUoVM9+7sazlbfl2ZdbOXv
I7u+lks8ys+kBkiRikO++xocvQ1I2L4m9D/8eBlYNx6y1zNlrdFMM8hyohRbJLa4cfrHqy7dtdMm
QLdz+LmhfNBd7+nUYhkkn5AK/Mif2lEzJvysmIfuXql4IJp6tYdLzr6aUmdvJu2qgUw073AeZlwN
xiEJUdmyzTrs2Qe1lIeGvrnltlpqZxNAwiRITZgCEtS6DpaJm9JMsbGO2bnu736VI56ArOFtlzCE
5pr4hmqKr1X9ki/sFdB1YXNuXXE8P4u4fcvytMRtJjzIns5EWnb7/E+6AX+lKyXT4/dmCAf5PYa4
1IiPC2N0Xrp4/ck6XWf5BUb3Y/wK8pMLexDCF+Z39lbKGT55i9fxSxLcLkssuSFFNvgPiXUd+Szq
D/y/0YR0OLd/4EDxkHkDYaKmqtBSdM3yIEZaTvjYC8Q0qyYhOWdFw7HaifTKaofqdPHIM4rRPnza
QSP1jjX+zyhrEuHLLh3f27cPdjaGa2x3j4BaeySmvoSlBbgQ9DguJtD4GPbLMvL+VGCMoGU4oaPs
+iWwq/h/jNQyP62psheZHEpmzxTAw76YVKYxNF2UsEJwbnjTrTZJHjBp/iNtjPby5W+BLRg0SSMn
Q06N9X3KzQ48Lg3VqUIvyJhotL4OopdaTeMDQexi/wq7k6zYO4vC5RgI7yYQddwhwd9K3faQC6bk
8nmylVDaLNiieR+vrWHBriIV3yUGhGZ1rF0X4uDyMno/Vc7M5O/MbaY63TS9YrtKQmc3q0t73Zel
xAS5co2PBLUqbBpW0anRVV2HdraCGla3tBNCYHSP4Vx/qmDBlKPvJDBI8PTztmY1HrLkSdA1W6eD
6eosAyHZIe9YfoSIi10tunAvEv5ChKlMafMB/DzWTQ2LlR8Sq8fWGeM/KAKNmvezhH9ngjG9++WN
ZhlxucgANDojR3MUXzD7IdAeMpB3aCK+ZZd1muHR6UrINmStRrbF8NzjsDfn1EJbDchS82QpAWeL
ht2REses50qOchSTj+zo6TYN6loQJtmpVMEoL9yNkfWoGfI7PT/iIwWVZXyhSlT/sRiZ7kTgkD/s
4OfAAjZPKFjlIOaQCCSWZhTnruYd4tvii+PJhADf5gaYf7OAjqRG3mwtuOlsXLeFOhpBu4euU2Mr
JRjs0hM6/9hl4xvfrwh7as6mrgSAQisuj28WS7PsX4FV5U3zwcnFSG76xMlQTKiNfCCFjpaXaows
BWkAn+SBJ+XskWlxTUe6ayy1ctWyu6qt2VcJW3rUYzv8EHJ7Yhkm4EnjEltH9TZZU0StemH/pA4+
xX1NNLoJe9OCSiY0RHknzk3jKZuOZFkvU5B7ieYQwuBPsu0L973eiXjNhcvvbsS6pdqlwcyaIoEC
jZSQcSobVifQ7qs9FZYqmIhkfDI62Hf6e0KJU/2+cPwcxgxnwB4WNdAS/9bXP6YJHX8ou57QflzZ
lShzamdEHx2Sb05LOFalNqTVQA+4da3wjPr01Ef2F4Vgcw3rUCcXbC2Ix2HxikFVpsYYrHZ3K3sY
undi60rF1mrFK2MMfiQ8/0dgmvnwsn3yLj7zZrWUYDS0UJhp3DgItkA76w2+ySRZbm8wuq/bEWl1
rTtzDzVkaRBRh5owuCSNxZQZhDkicBTkuzcFRFe9DBiUDWcnY0FqeuHPCAtPjqrOYhWUClsbpxoJ
LYf/wMsO304BXBWvesEGAx0FpqTLBxQEZTnuoNddOgpf6xqKpjkFOUtiQ6tKJNgRQHPb0B8afGtl
cLXFLY8fGVFq0Rg7xiWUN9F3cXQgS0hPWnK8nerGct1SdAf/W3tYB9YllDIrkAyXvKS46h38Be3D
dX1NJ3m+6s/bkqmGgADYzh3aVTqZkCva+Ib2RnSRIXVcLFuvPFChJ4IYM72yIWMDpGSAkZOr3W3X
WnBjyOLdliDbz1lNsVJZbUF8S7QS8Kox4F3f5D/o/OIZc4c+H/efiudbp0L42ijGa1D36VDKhf5e
gLyXhnlTI90dMjXeEv2FtpiiO4rbjY3Cvl0b/DtjTVfIilP5SA4YXBvTWCLyYQo/f8Xauw+UCMQ/
kv+MyVJQbhuUh3aC1/slZCktC4/ga7UVqP9riTL/P7VIs0dBK1RyFaX6m7rYgvJ2Do4Lo81foaKU
winbOlYghRQeP6xQQCkvsjCcLB2auLxQM5fdGo3eC2WTSBfGsbchntaXTWTlbq7+80Tq6tcVC/FA
aSIYlkaC1NozW3N5BZzJjwag6e7+MMTMjWAkCjxJUAErYgec8J+SsielAeCXO1T0hD1ymfIrp01+
CWAlxNJUwH0dyGIKGLFpoyLfB7+NZhijeNwxmlvAkBTNJKzfYuUL8fbI9iNIJKt093SAdumv0ObC
WiEvVbQXKRAxQxjldyKfXmSUdgJ5MEFkVULO9YO7zY2uc7lxIZmf8hMTpTXxr2QAL/pIL9ZAbruJ
bbaTtar8WWebTtx8ZnAxY+mmyyOdklgUv8sgfmwwUShQrgjVBwqm0Po3+vEq4I7hfBsEufMO/8+1
DAyg6n7KRhGteE0ebVPKYjKcdunP3CggToMQ0ctV+iXs/2LWdmfaW93mfFvsqazdfI2q1xZKiE6j
PjV+IiuZfxJWzDvB1POGuZgNho5moG7jEod0pWfnJxfJTY7PADU2e3n4KaWUpse0E2ZCHOtPxfZ1
EjKYzSWQMX+4i8WDPhLuJGhPLvp7Wj2sNejmNdI6+mEkzXY1JMF0ZHiwMhFvIipLFsViBVC5UQ1v
vg2NrAM3Kbdc76RTiQjjt7I6SO+QGM25eFgnDFXlT20DiFvuGwVwzhF2aCkgDAbOb2iVfWLySrgT
lO/J2j5MfE724uepql/LtopbcOZkuRwRpHbj4HsRvntVQ7N7ErXH280Kixuq4NodnCbj+2kFP/G8
JdmPYwakrbCry6g/bPiqE32DWXFRDTyI0kMygLarnWH2/ZbtCd5gwQLR/nRFqmH29x//B+KXu3o7
Mn0unXfqDUT2Da+Z/BVWAW6zEkprIartE+xqnwzu3qB93rol2cbma+A+kAcsn/oaW03coZTfBkvt
fAfAeWY1bk3qhPUTf81rUR2ZiPxrTAQLQklbcow5XFc1ehEo6Av4LKSfEQUGtooGo6+MTd7zgXOp
irnuD1gK367ck1imr/MVR9hALPN4ysBT2KVT8uPFBwb/jGVhvZLInCkASVUPXTbKZcslA0kU4IdT
Jnb04A/vLAElfEHwvKBkAXeRw00mvclZVjMOYm41Lu3aw4z1s/yKi3hiUamjtLGQ80Vrppm4+np3
PzgcYnrAy786NgkfLA0SyPgIlLT5B345tcCp3K15T7Pz2jtP9I9BY//TcdqpzFRXz1FOqIVKxZ3Z
B8xR3oRhI3i+MJNz5ZX0rcufUBHPsgzHh1luLkD1O+7genenlvkVAdg5qabc7JRlpCBPXug6L8R4
abG46uHKEG9VB5U6HxFrN8SEXL1/lxHg/wUCJoLsjs0F3FmQkAtbmUv+5g5wFVLc2Id2ME0lUa1y
7Fa4nTjSTl8wmqB1XMi9u0xnUfewP4I+LZFLMrHuWbw3LyoEaVQQsfGniK8W+XvBWTKrAzOQHZR0
c+kWw8osbAQ0cQZgwCYLoddp+0ANIpGjxZ58rRgZaCq6QsglkbEyagds2yfNg1vetbdUDRptvPAM
FYvJcRvywscf+5oyBc0CcLzlOCuimLjqXA89ifmeDYl6YZwd1ioUp407WI/XC9+rvkkU+JjZwFrp
2A6KPONQ3568yP+PUHaXOfz1cxXP1h1QI8XLEZgU8CAChLVJfwb6gF6Fr+xuhDJCBHlKiJ8Mm51j
2YDXiCFl7IMyzaUa248HR3WKYsKg/cZO/e3iL1NudchIBgtXiCeuNT5BaWp4hVMwLho3s0nHRP61
iZ0P2xG/YdzMftk8mJ8CrynzsAXXTlUinKs3Q+CqNr1yRk62mapOm79lE0xx35E0chlXW6gyoOTn
vobv5gFgEu8noqL+Inwr6e5ViFWoR6z5xEjAtUI1SWEm4dFKk9lvVP7zE7RGlTFUCfs46ZPIH5H2
3qWUoeETA/PIW79eEq2Ep8e+ejE+FrN7nh4QAO3l8dETeuZOZx5Rtjo+zjaTbyhbP0eYv951cNxe
UxqvcmoMRxafMJFpLtw8sb023ME0jA/U82xgOmioC/LwgskdWTIuKH9Z1rGlKzmDNHJFg6mxjpNP
q3pY8oZ8/HpL8bpJhNeK4kU71kInF9zY1ThR7YGdOdoDg4LzEtSPeoNzK+gnmjjOVQTGkRw+bW28
U4xCbFIjdiytVwN1gICWgTiZfc7c2OHoQ41Nw0Y8cTioYAeAY90LIMD49gpvV4pphorBbga+LMoc
QypKlFHo1VAUg2wgjhPEeBUQ5F1uQ3aTcLhNRP4TjCwz3xy632DAxJgIZgZJYIqdlnVemEqZl5cb
z2G2TQF8Lkzh25G75hQpkTx8UeLJ66XsXLXG9rstR8Gn5un53e6otPWEIaGG+XqxVDyUggz5++Wh
JPl2TjmRjfXKgvOMigaCvaOtk8EK7vJSmHA1a3KPiYXzk73ViF8OXl51nCfMXXmYT+Rbu1O4L4mP
UuF6ZttSaJNrtWadeNOGl5+eMtRmMrMc203PWn6eltOf05uh8N5LZfmaCw3e1ovUsLscEIlHeU2k
Hs0SjWf9/GMWXTXmzQUaOFPrlm5Q/a0YiG5C2cvJmNcFzav5gGF31J2GOgoGh6a/l4HYbf709q1l
txXa9SybBAYtL6nqvAjpkOR5yYQuvpYB9JKzBdTkGh4bhAIejWqwQK6Yk/J7d/ylrMRmKKb9l5Ei
M++rKpb0cuUguzvT2XhxHL81baPKUrULS6cZRZwvdkPNBZPHmkbtkSha1QgDvP3szOycRRxGuA58
K7848kBSmXrowAw6f1ESWVF59Gf0IefUlMpfZ76aRQY3fvcrOGU/gaqW2naGbdTftd4Xw2ZxSwoW
4978uDTG/cO6GukIgpDGxn79E8SGcc2mV8zp7aV+CqD8SalNFLrcatKICrPlAM3OpBigM6MVX95i
T6G16ZG1V5iw3g6g2jWwpxCo3+HyZ5up6fcvMlmuFdNBbgGNPKNR/ujaf5jWVsPFeXc+GafAxiVR
3N0RiRbrXQSXQcWbzb7nnRz86z/vVf5CjuivKKrIe8OMMQHj38HvLyGcZ47vvHdd+gAZ77eaFW7L
/bCborOkrsOTDQNhaB69CuqKQ3te+XQZoGIVROa5PoCr7UYIvz/k56aLZs6HdsHnW189FQ2TUcwB
p3FoOglZSRRcZhz1MlCYGyJfhWoY/kEpYzIT0JEoVXnyCyd7gw50ZBPlGXdrc4ZVPBJ4HKb5RPwJ
QNSDQPOsULMGrKr8o/psbgI2J2MB/lmLC1Qs/phvF7DjXzle4VDsfs/9eduHYTE+hjoddAOQf/hP
IxbhsB1yMw2LfIEznlPwS916YsrqGBhi/RrzrwVXc1OfS0ZXvBFD4pTDRK5KzAcTxxKKVcs1c3by
k9UdvYUyNoEFzF3YKRHtmYxiyOTi16rVVXzfQkD4pxr7Q9vRZeEjYVccUfklnjOpN6i/tJmDizXW
i/OMAziqNcIymlh5R5fjYKAyc/wRMIhf9reF1xRBUjuMGmhr+qAL25rOEIUzlFIsJxBU8ifV6EfT
yrr3APHymloRRGPx3FZmCPHLlYXuKeCAyZDVbStWW49Sgh97GYSeoB0ChQgo33jTtIznAsgWzW53
tMbWhkx3t5sehmTHJ7P1Ak8S+VKW/mNW5CFO0SQcrcz2PssK7cWQqfqkGqZDROhUlChn0dvNfpif
rES4WETflUZKn5WCZeJE6lY3NYLcheJ8l5NFN9W4RgADVPY4zftxxIhpE84zrT7MwZJDrlxL+064
S+EJUk0FIcywM5Ra0XQs5bEsetfQeJjKjEJaDs6GfgA7JOrj9yDj5oHvx0RLZ92tHQFDzbiTU/WA
hB+iZirAQXqNkje80VJiWMWBcnvxWsiVoeAl2C/KO8abIEWP8cNmXqYs1vgvWBIeoTbuAWXp7jhV
MlmTF+6QvKJD1OXFUKABbW65XJIF17hx31HWYM6pcWb6KJ/J/ZOFlChoX2q9GVjPiKTi5BSrlU5R
ySyZ093KtzlnZkdKV1LQU9spPD7NyyNqw+tZXcF5G8YjRClLiXIE5f1tnICj75fxhmbQN+VGjPj5
VAXAXAbct6VG/61F1SwEDbFqtMdFjI8xvXjct6J+iG8xwkc/cBBJF2E4Gj+v47q8FugB4RX2f4g4
ze+Od2HFOlOVg0vYIaNVezmL/Yy8fJkKn4ttn9pJJ4hY5B057ObrWrnN/aBMWrLhWSInm7ur7Rdo
VhfoImZwtYzO9uLsTfdGCu0OzlpNlH8q55QXZe/rQKa+PD85aw4hcr8R5Wc+MK+7u+7+oi8LjDBb
1+RbM9c84tNuWzUM/D3Lp4l2XnP6R1sSUNQKvgLp+h1ZLKqRqavJ+2kA34s5dRLTW+xNo+tJz0Hm
PzaaBEhXclEsIEBRFhoyBMGGyINEW/GnKt+ZKtXgYykn49AhpKfMPWle3LlWzzX+yumqiS0Hz7aq
g4jHlcTH6SJKqyF3QCSGulJRykVAb3L7wAqlR+bU+pcPZwv73EJgL5YYU9Di5Y888UqGE340J/ZZ
/i1BMRmN9zUozgmAYSLhNbj0XXZWm3zgVw4xOgZ+BwuX2P1OHjjkedJHaiFy4FD9MInXckiWDrbo
1IPjkiQ/RKp410adkjxGq7WqRIx0MbgY/idRBQc45CeuXZL1f+uSQBBnuXXTzo4rLrAL5HNmXomL
Ry6IqrRqRdIkTmE2Rhkrv0vHIBYxzI5cp23AMNX4SAgrEIwXM5k1CM3wtyPNR8ckgYr3p90tVSio
YPavA2cvZtiyklIz14IK12f5UioA+6Mk6u3Ud8+NlRxfeLnWh7JOF/laVc9eZiGQkL9oJ3YpD3+4
gkFJunn+W7oOlyZwSEruSg+CpasuxXQXgL1MvnHa/+jECD6rbfG+0aSY1pBrA/hzfHUeox2YKj2o
y8QVVIVu/WRy77wyp/k8srxjMVzEtfdLq6tnQqvk/UFgO1rp9nkoW9nQTMHqNso7PnYr/8g0yvDx
IM3nIylYb4G5lajk7EHInnKc2U5ePivVab4JUMsXMzqY78R2jBIqB3ZaCED5Gtn2B7+oJ1mUOIWX
75zjSpgXcnSVTmt5oqAMkzUWyDdquvCVKBoYuTgo09MFmoLkqxm7Xqf7Y3toQ6FEfyQb2BXPL4wH
XIcKMu7yLcPkU8XLCvLqE4TZBQ02IbjTaqWw529PviRhMaXV8MzCnrRaNsd0nPD2huD3s+sMKoNz
lv43pKZG3FdbefhHwEG3trZKGr5KKUJ8ch5nNmkm44vzCqsZJIlquKjgWQJ3MjtL3rFMirDdeWYj
orPGHhcQe8xGVVwGJ2nyXYBT84fJpHT/U8tFmaer+JKq/U5/n7FBLNyoHuKmSiaxZUo6oc9A9v3G
LCv2Iwx2WAAY4BNUY55/3fzouwL80Flt4iafHsUiIo2GSZoQYA4RBj/iZ8P79ppPsf6o7TSPHX7A
ekz9kn9dpBNpQ3PbAO61+LuHI/KpSyHLFz2k9S18Nx7llDHBPphUutgcTtMV1u/RodsTmD6i0xZK
7hjS7mLe0KxqmdNmB90NVW3vzA3FxZnJvpaLh4ERm6yLaRM6Ux4ESEOOWiupsj0qtGJzdH0OQEni
qdhwIFqXJxAjKxYmocCDZO9YcjCPt+LAQblr8pKZHeq3e2ZE0QUrwSVeLEJgOx+5j0+LPcD0Ssnb
UFSq4wDvhTSgejDv15+QrWllcRCGbGMXx8XnXJDlhXaSBFslAL/TVxW8kJU7Tl09m7Y5UnvX7DQZ
4bnJh8MeXBv3VBc3U7teT7HNR821dG/MtJYujdwpRS351XqzjGGPLnVJdQu0tikT3WCURD+S8wGk
4Ji4UxvkD0a1Fb+twWyuMOSEH4ewDLCuotEVIOxVANJEKhCS158PzRgQU+rovoJ82Z3Eb15Kjjjk
gc7pdvldRO+zqm3f2/25qfgkzqQzorPDvfsYCdF23Oh9Gy5qnEbV3wyoWCg+BQ3tzo2YHphn1dyG
5KBnkYXpL4c+cAulQOsc+2AuR1ADp54SSgABi9PZzDMSx2eG/B8uMQG9Qoc1Uuobkz5B2aHNMvEt
tXTBXSYak2nUf2vsi8J68D6FUi/0idBShzTB8keL8aOgAHz9R/jVPHgYDyviPVx2rceaMBP4tsx0
nVh57BNJREo1NLCsTgLP+mrS7/vS5DxrFPQo38o3UykUMuw54+rzP3t4qMlEy8P1c1h2D19TT9ON
9eIM4LRDg2h8+n64XQywsJ+ApWPA35eSzMpW1AUYfPr7+Xl5DFOIyAyj7AG+KN7GBAheHexbuM/V
p5LPlujqDXiR8QX2ghBBcut6+cggNdfRjwmUNBAO8D/Rnp5tqlA7qr7TK/NttShGeZvuQkpgnMiY
NCEFR+RPSy2tj5FZr2WnSX5watsAObYaDx2zcXd05GPV7fQiMuHqn38GY7FHWBobhovQBbVzrZtS
I5IEFeGUYtj/YrUhGCsTAaPXqOEpu8HiiyiPkZreBK8/kGvGrK7CiGKqlzGgFYh3gLzszLqHswur
wKolWFMRHtYq2GJFMXdWljGhouh9KH8Pm2D6spsN9crS8g25YDxzRHM4zmzaiAFAoP08j9s7sP/1
+aHrKu6eZ1eJTNGj2nhkLWrnoRil1RmaFeKZyWJptGdVAR9fV/kKU95JziGenehqcVblBBXaVCEB
OGHQ1XSRUyDbKDU/vRFNWXOfRMMq05YOasboH1hxsRv0yD+wcDmKJn4zLJ3/MnRsVRlJnTe69e3A
molmDBtmNAX8ZACdRDpyRKtqNiKrgS5cQusZ3zUpryTLY4TY+iEBPRFOPjoCevjJFz+QAR4nvrPr
AfTln5WX/hOx9/bZwOmrKv7ePN64TI0J40H1jaKiMPrWCk95hP84OZrIQlt/43zasawM4g38JJZn
U80hcxtPgupJPkn0HQFijV8v3+KAwZHP/ZyAjTHjK09aIJAUx07XBtOZ7qCNfounWPNTBbyPIJ0p
CMjH/HluCXoStlWyDbfJmlAx67M848leI3mKxUw8+0Kqd7PhvmURQIBuxEg0dKDwWuaAFBhIYua6
zGzBW1IeXNuP3o/uoqgh18T2uTXLuqsPTy3Dv8nQktWIqllI+qKkZNrk6q2XnByG9iyco4RGvdPh
8DXvgYPFd6eGUn2uDtZ2BQjs4V9jdngtQA6aYEFwi4qBE5WbRJwTAkgEZVumRRyc5t5JEVCw7PyN
ALp1U33xg3f6kWrm/Ew9zNXgtJe0uRjKHwq7fcEzg/11hmfdppoX18PGBe7sDgRqmdCbhk0VEjHg
M4ltbD1+kSlifT1jcXdpEVT/I9ucxJjv4ucvd+nAlZ791s4Lq8FY90832tHzcm3xLTgMceSo/Zn6
FwZ6K6EYepMoTRTjniewApDIZVQemMED9RqMKQxTlKIUuelu27/LR87gXl+GVA09E73o19n4jnJH
E3UgA3ccyOLGJ8qOGEsZmjmGI7wgKrIlSt+gOjE2e9uO5KNtH2HaXLkouEjvTb6AQUV30vOJhREr
TPb9dpt8gfZJN2SPEdd5JrXGUCmjqV3yhYMdqdkR9EciQy3CovFG+lM5bsrd4tM9zw+coQs+/0ab
pap3wKiSBZ2NdJ4heWbNoVxsTQUl0eBbB3TSSxm4eGzT7Rpv4RMvyAVVdIj/CalPWRskdViyfG5p
orHnjqctz6Zgr0HmPRcpbCXrYxLlYEmMbmN9Mmwy84Be785FdLt0rxEvDpoQdWswyq6JsQmZ0ijC
51zpmSTnyVIUWd+QLcgqnD0BUZ2ulr2pygapvVo0Q7XKKQNxPK9/XNDGAnhpYzv7GsX6c4TsHbHL
nsyFmf4nsD+ICpPAGrZGkS/fp6PF8/M9G6lH4xsGSBJsOihrKtK9kRUjFXCFjpMe/z0icrdChR6e
NRX/oWZo655qCdM/Z863Y/ENhOB9T1lVfLcdlJsU0lkKt2m5PejYJpX3s3vWJkerZYCgJCmtcbkR
DqyQ+PJ6CCU7Rva55CY/ajg0NgCjkgUlpoe3x5gAxz6NlgUgLouExegfR0+o95szTl2Ohg9UGved
5GmCglLZO8fvWqIXlT4PdxS8+OFWQuuWZFHV/Ptpha5fY1vpVzp7IdKHc5PWErO1zw5WIvscnQoD
+yfXH4szpn8MU+B5GcpeLAc8h7Ga6yVGvxpkkcXE/DLOVm21bdnuL5TdkX78RPcUrnSiasmWPghi
4YQRizHoYKmzIn+LYR8s9jrhZVv6nLWWwn9zcHsC+WoU+gd5ImCQSeqX2lfNL9QFvkWY8vs/BKvb
sAAmh8HfYI+Ixv7nG1af5E9DTV9FD6lmpg06YC1ySYlxTtNIWXQyMIQxXOf1FWN2czl4+WDR+AXQ
c/9stN2EktDHzaLyh7McJPcYIF0LFqk2fja9ZwKzyHZ/vGTMwu2XpMam7SP30a/d4hmzEFjZ09ny
FMNOLzaNWSrsaFS4sYbOQz9uB3FsYndB0iwfpOlWeylWZuHUR4ecgrarT9lHRG67zxkruX0mWeiq
f5RlOTj7K0dtsZ3xOcpt+voqVBIuQC2yRtMi7fCwTu9+go0EW89qA6pVuRYGdc+hE9gbAgl3uz75
zdwTF8t9lhhbBShKAQMMiDIuiKn2Q+xL9Ovv4IhW1hMp2APBAn2rVYaPw00yBjpYGFGNGC+gYie8
nQ+i38obx5UOIqGOK+7HE5mZy60DXc5aJJYIctEPqM8rAtpibFS0MjhKMOQmx36oR1Dpf3+4rq5h
HZmwy3AeV2m1B0dyx8iLScKhVqW5qOyT/hmGypGhVvt/beGIeH276vpZmwBrwab7Wn4gqleLWjdp
00rtu4M3oaVsJBf/vDJ5bCbVmvLpyd8r0OAXWLIfOPfjfDtsKtz8cPShnC1h7OEZLdXigkwxIBuV
SgpYWXyuEmjfNxATqMvPtLNWhGgHiMRvR8fr6rq+FF7LWgV4cKKwBNFbOLsiKVROEzCc6fXFg0yH
e+MXXiTO//ges+32ebuHrbdzhn3n+9Ifvrngs8hPOPfIXFjkBxMdEwdtvV9RFIVvo2d88CWhe8Lc
KX39xUkbWQPe1VDpYtoAy4MZu906fIjbRFhyz+qKR9DlmoXD70+32ZYkhuWFXnbbSHr1LMb56ED0
hUCu87nbyQu7Ie0+jASK4R9REekuOpMVC4Va/Cp/4AkQmyytgrkgX41EDrsx+7EuJvslL2krHAtt
7SJ3jtZq6uWxrHhgkF+q70cUb7Q7XHZIpuKYLDVLeQZBdDpVRL7YFS9SPS+wJ2m0u4taya6Cu0Jn
f5VXc919FJcULXUbyH4XQ+GDOQ1QaWJOoiEyzpxRnqiHonM+7zQeTm//b4j9cDeYFNXTbcz8WP5D
g3NytYhMBaT7S1Zk8OIXK0gOTDxKDQOqZAEV5wdj0uYpHCXu7b5bl0ot9LthN3oMqndjhqmhQXHf
t8yn8cJ0CYRQiC7nIAzQjxnA+h02NAFnx9l6YUskZUGKnvQJfv/DyMnqR8t4t28qn0hR5C2rTrpF
e7DxGLRnBxhM5Cp008iP1+r9z+8ULUy7OzrtBknyXFzeEy0JxG7xwQDW1DOr48BG37uS+2ttTnhM
MFt3biJmEe7nmBJDZy+w9oveOQsR9k1Li6KJV0+HvLkpHvOTMPmcW3BgwKWi06g66yyD7r9zV24H
FsCLgXKYzVTpGrovCZO4J2yo5VHbl1dDkNj7mZUQSX3yeH0HdmQcZ+p0ds0bapGf/f4AujDCGVDO
LjHDfZrfOuicYHR6A5LVJHsjJqiMhqG2MHdIyo8kHrFHiX2ZVd19JjKfJ/gSCEd74ojC2MwMbC7D
iupAQrFW1QaztF4EfGI0OOz0S2/LYR1oAqdgcgaJ9D7+vfkuWTcv3ttDe9qzULysO14KccnNGg89
FTQYb7HFPOxqkUlamsU5SAs1XIMSqjEQexdfOEj1A3LEyLE7I2JZUi/mhiAxVSEd6xsf4kJ4O15j
XEj6N++uHqZiU+0oONzh+vZIFKEPNw0+ssB1VoNxYoytL+QjsRnou/q04wHcaaJ69rkJK08D4p2N
Qgn/WmM5grh10QoJmvtbuxUfs8jHBiuKAaazKv1kAEo+SEBseO9cZ8+MlRWsxh5xubfodfGAwtnO
1Xc/loVGYwSonzpKVPDWe5LQkX/lfJf7rLTLhnqgX8aHjmEtkF/J4q11FFv5L/9djqhK/w+NExO5
ibpoko1qJU+40CcK9bPOGzer+BuFb2W4elC1ARNc6fUXWSVIiaVPnRJO1gFtkjHMVksgbGM4tX8s
xJjAxhVcPkUQwYwJvzHkxr1Edp/eAxCiLpEWXOGCSXmo5z1n50aTFGU6DgMc/JuMolDTFPQs8qH/
HVhXcKyujvWM055PPNSKx4Y0ZB4nNsCH4caQexd/r8w11jHmxWnZCTLv0snQv4onXuPxK1WUn0Gn
7s8W7dnc22w+gYzAlpmSM1SvXeGvYIOofikHH+3FYeBJfKGlaSiiZTccHcURyEZZ2JRC2itU5BEA
A5a4e+RdRkLX2EH707YBL0QEvjUokmycizl8jEus0ZMcO1KelI21ppIPqffXH7LZI3SzewfM8nhe
jF/U4MK3DJhaXiPEmy1Viz5FAFG8o4HHDzhZ0v+dkz+wS+ucB6idGsT/rjz/1BP/MFFj0CelSs5j
olkjW1+OcvHdEhjHn/z1pnOqXlcDVnqjkP/kjW7sQpXVUEtpKOQGyBK9k3zPzXWlJyCvloc3+KXp
ECCLteoEpoMVCysSxkwOGTvcXS7ZIF45wr25Gy9sgEOxR5rvOEKsq7ULXLUH0st8eDa9Ekfpt9zI
YzdgW7e1KsDCHek+PUmPSweXZT7eMyWaCAOZw7qQgsUjr6Fx91htUO8IEIK0APlhFm4zezIouZDu
vNfbOgYw7bdUEVtPLhkjJUz/b0Z5uBZK1pTsjktITT1+5Dg+n9z5aLobAoZwdoSDJXkCfE4ZEz6C
pzW4AaS6uwf91wEAxIIW3qoqk6Gqw4JjZ3y4sWMp+6/e/fJ1KD5cLMWquCD7aZUq1a1uapsTFDcc
dlgeoccaAkogdMF6UJ5I7E99QiWzwqlpJJeL7oxpVIufHE+gt4NQFWyQY0mD8JwHUXc6HxpTiH6H
jwqApqLa0/om8Zf7SvjMuuiL0Kk6K6FLSLs/a4EXu+Pz0lGpCNGPtDCyDWfdJDkY5wjTvnc7FA+U
V+JZAjgW2jXUB5hsaFgF39xRhkpE2tK4EXZPk774lcgCmKRcTWoV5VdcfdMAgXF/WYP6WiJn+G4x
MD2r3AyHAkxfDEU/MIaa9+HwCAts60tJBUcUW/d/wAdY0VoSgxzc283PTawH4Le5c1Z9yxMMUiFD
J5ujjvxt2vKlfQxbNKv3QSc7WVJzJMw+FsU829DUvT/KahSkKlKOT39N7hYzYQjVJoMfZLSdGu2Z
N1XmuSB67vFxfpF8X4UKgRwS9NRH5qbsYSc0O4GmSB/jPvmb5jUDVtFlkctY/FBvBPOec5ILwraQ
tcPnNCkK7GxxMbsiBBDO8IlcJnA7iPUN8fLWr5uN7nKq3NP4i/xnkxEFXiOohH4uiF2WhmOrqCGC
t9vTSFegxMladjiIJqitNzoAD9j7u7wXQ0KQHZTkeHS91XwQ4qjxUsE73aKpw4juYyg1ImYPchCX
w5CkaoVtO4hYG3KoXJolW7waHbQgymUdIxtrOdADjuFT6vmtBmleVw==
`pragma protect end_protected
