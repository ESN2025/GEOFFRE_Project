// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:26:07 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YzyX31LT1wJa6UN3+GX8qZrO9LdJ1oNgT69XLGmQc7sSgFDsJNuSl/uH7pH0gfxx
dkusAgliJhmc7z++Xhf8whONw2D0LgIlXYYMKfTmBpU4PCOpI1yvJmBxydNsBIoK
6rau2WMM47NZzXMWrB3ugIEiWYBRhuT01cnA/B3LvLE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 39552)
2derVBz9IJ4qHAnk/+9grGTqAZvsKQ+nmBwSZxzDRQY+o02s3UdwpLiaSJa5xjh2
kEpxBrGXXTX4ghntC/6QRTSTUXGSGrylZ+kF/flwoj/l2KHAdr/Qk6v5K0TgAVsA
EaV1/rfot4uqg+YhPnzWo9Dp3gKbz+Qr0iJ8jBXi0mCF+AZJKDiklZlFF5q1Txx6
nf40Os1flV9qcsCuplQ/pHfPwYWHvRDQQHGoENW8NGo4ojD2jhO2awfAvsOj0jYH
ziOZGajLFsQVDDzp1BI9O8aYnsxSfTCzxlxmVnReYW7SFDXy+sLdnzvJoXMHCpTr
+zjNuF9V4o0LHScblwp8KLve3dURlgu1qDUNZUU+qBbwQyK05j8NDbaxx+Rpdj7H
A/QeS1FilbgYnHSRs982nCNNq7mhuHNZp25PqfoKHoQa1JQRH4Rsdxyrhjv3+Z8d
onid34FyKNkR3bGs8x1BgAiyKbnEUZV66vcXUR58OS95N02nPR7AuPJ88X6Sj4Y2
BjKrd6o5eqc7Z+BN0tbrd5esNBDkrrcb1IITPr9lutEAw9iwVGwX7KJbH/E5gkLF
FhhYDsXAcMuskKdSe5jE/ub1x4QmY4h+ZfIuG6oYlbx6jn19Q22go/6XhT8q+T1R
jnWLGO3VpCBaM/t9+m4kHgqiYommgLXLB2wdftHw/ePKDbeKneiGSKSxy5qTYfle
Nxlv82h1UyInfmyLXVwl4TGLMg3qQ42cZjyFZUKdce4lQ9QkBbJV+LMWcUTkDNVd
aQUJYsh+SOTn8aRQWtpy9XKhe2GMyVrOa2H0EwrOIl9Vk7LMX5Ob2Mk/00i2YxwS
0j7r7YPwXA1C0cBoAZohcWrCQOoAdHjhES6RqEant4DEguwX0dG/SUJKqfeI6XbC
m6BvcBXqRRWk0vVOh1Sd1vwskyHOGsvS7KjCjNfqmEYU32ob+OgTobyiCV/dN/Dv
sEwSgQudNSjAP2ux0iQEsOPrtoaXyHA7PvsDdKPBb3HWmqtIzXhBGKbvlSw0c6U4
kkY6ZZIXjp61HmjQWftxLXLNIM2BHKGpb1K4bRnpS0kH3zo1bENMIobpWjxSMqYn
sLF52/JTuZHGTRPIulFzPO53Vq7aM/yGhI0lvvnJPeOP7hAYJx8iNQP0eaxYkcV1
9S7K53F7Y7YoOknuePHb4qUyETwHmxnBnevNZrkt7ESEhGIM5dq+vPzYTJJKH/Et
UaINThnFshJB1g1GacQDoDjYXdhHiFZL69mwEUglg8NZ/xIDgQY9ZmUZ4tvlDM59
MAKxiqAp8qIZmSEjqWPEO//6pVEk6rjNfAkpy1Y3QNTlT4WnNNZ/epvmkeFq0hQo
8BUo03WajOS49OENLlM3hVbtbT9CrD37gRNxfkeXxB0NiUnDicI0Lur4SedeBsxS
ENR1qDOi+iIwLI2dynAZDQxD7oDRPJX/q7trFYQi+Nom6RhF8PvMh/fkv4wiadBh
BfuYWYYmr4i6hKjG12OFhw1hAx29ZnFAKIKtwY5UT/okroCQaB/C8qQ+vky/m93u
TsRwrpnNaAo4E9uuZjj5rjQRU90as307q7Ww173/TY8hNZGijLxstDyeZyfu0LXr
YCQch27W/dEY5LQXnztbgMnozp8N0sGQrgpnc8G2r8pfwD2V+4vC0vA2pE5YLFVL
yf95W94dgKbpsjYDnphUEtlBor9ekh1m+gddeiU41K5DrQcWmPpF71d2vi/KI+QU
1c7d7wB7cC/pNxht53/7Lw43a1DucYHjWIzBfY9LZc41RtJi71Msvs11EVZdOd/d
RwMg2AaJtNRYAqQpi3z3JqDdCNxRjKkhQLVlL4BkwHCc9KVNc/7ETB7lEw4rduRA
y3AO4qC2m7qjQ8jhobbd3l2VMvVBIBl3J8fm4tjQ+FT6HU7BFGZojdseIqZ6rorz
/ulvPnGbBbYa5OePUOkTZxTXsl7V1aoCAxkNyZJTzEdjrSbZ1SAjnGQEJctTbyWZ
BlZPVMZFea+X2CePLcC6mmn7YHB6XDuUtSiXC9kEoPHMh/ZrjO5bv8lhgjMMIdDj
vpXsBCQZQutBcodk3AxdP55rNHCEKhuFwMHX4GQDkylsrV2rT1FegpgLIKp36IML
3UeOu4rP0NvaW+Ja+M4VsqSQzXF6FOhzydsTD09esFKSONDGn0ewsvH7C4pyfasF
q8C/9d2mJDxoaXFIxARtEE5WRrXDmlHLUuCV3akPR/58dhIPGKRtrqHhWF49dClr
tbDcCaevvTlrB/3pxRWtI+yh5K6v7qtbw+0FAFWyXrs32ZGj6AuQ3TYqtP8tfCq5
oFTW7dvfP7DO2XI1AH/GNLbRi7NKrpHdYDqiCh6bdp/EU8uin+H95uuEtwH9aIeL
Q+LzAyegkOxTiUIE41LLPUxce9EruV2fMPWps7LyowVAS4ufPGT1GOWC4wK740tV
tlxnpKsAk0M0hVQznyAQKa1zpHeyHhEnzrzhy2HG2gZuuH3mtY7ewtVGVkGpbxOE
OeI5xUpril5wvO0oOJnyfsDESp7vCFI/812gwZtxOTRLuTIvBdG5WrjngzTSF9yk
+XVCZtIDbwTJPa0C+4oAC7UkixuBDie4lTz0K60gHyV1i9z9XJm0QhVQzf2it1yd
LnHANGYsRvMUio97A89D0r6F93y+NV2qgMVWELTCwXf+20PbCIkRIfzc4VsfmE/N
cBbwizkmozqtSdF1VhpL7UfELbY4Lpm/ndyjwZE58UuROiiNl767idE6aaTZavnO
3y/OBSLB5g8i6HFF6dnmosryPc2xPdIkjzDWvGTnHatxgjJwlukWOUMeyTYomGzt
7lMPmPDJCXFGxG1bkt1JaoHaPa6iRxyU2uGuOfOmWjHkjwUoy0w7rEqMBeiwdfG2
vDGq8qF7DKClDJDozF52tGRVrhwFG7dO+6/bQhDBoIW59JQExGoF5rLvCr/X2NNS
3NCnH7QQTihSPG/dnptsVV1Hpe8yKJYgAPvdKFmD70cCy5WXszSUygHF2X1aqwGB
5JXD1Olay48UjFUEO0VKA+kUU/ptLQSxAD8VJXTnP4WDrBXZAcBmvRWyalMghthP
V1UHt3Mghp+PSMuKzQd8mHfd7rCPBqHTKOI4k4uHHUAhjttUQlhP5bbTfpcS3LE8
kY8fFQutIGXyCQ0E/C0bYMHk14KLdOhhrC1ZwX38kAsBud0dvrP8Cr1GtJC5ue++
BYgDRauDUamaz0UpffiznsksBiq6cioX3icbdCL81bIHzSGbr7sIrTF/C05Zl0A1
Zzf3KQeIqAlipo8q4X5SjfSt7naP8AjofEJn2JClnnrPI+glqTKvDEb1WVbyhD/5
IDFLTuRNMc7QhrdJz+PAPtVQB4zJCdkPHUrLaB+uLlU7sOx6cHrPDdC8RD8hEeLh
nNyC06iXtyNdVDs7zfQwzWDdXM47TopW/DKM2mU+sFTNBK5FOtQbBGTLUKU+vlDF
FOKaswsuYKznuXLrGwV7sBbD+7QTESmEzdQh0KfuzAOaAwSH6uyAwD0nh+h6LAtV
3ZSXJzDPb7teWgzPgT9/5DQ2jCgaTyJNyTv4SX9ZwEiw4Ot6ZoiVaYEE4TtfVXCL
oCXzIFsxoBDwkcEdWqVV8udpEau69TsGD7bfwOAqs3Owc2AIqlNFpakb7Krx5tOc
vYdG8NNfFucs82Npraje3a+hGUOPdsKq0zgaTDG7Xgl3EtNSQCxe6yyTfdI2Fwoy
DfA8QdJeZ0oZu+WOqtdVayc89h45Q+YAT4VKZKodKj99phnXo/1CVZU9fMIBFd/D
WbFBJxgyYthXiQ1lD+YOqEMJ57uDXwU8Y5uEAXHn81wrVO8Qsio60rvTQ97EkVjC
LE60KnH/GryscuSimxOjcK6qa/2y3BIJjkHn23K6xA9HgbTiBDY3SqWKXpIER2XK
2wTGpSQR0MSpsBM5WvQblur4z1llZiWrglw2B+mfqYWKgx0M+gUTdnbEvl8VHYNF
ZNwPalQxapxI4wnN3evsRairhEBdwl4/fZw8W7ExAmWL+JGLMVho4g7ycqMiAqhJ
k+5rlsck03hETQz94OltWdwxQ3XZPrclaPqrSGY665tTU62a11TZIb0APP8sK4wJ
2LDr1skcjCHPWaYfEgx++JZw4LPGypIf0xmTToFhCr4RQUdDMfPrM/cjbCtnFSwj
kEEDCQQN5dtCfXycq/I6M6BK/qcAkZmz3k7egSiaY9AmdrwZT97y8oOsXfFHyzaT
6/VonITwlFVis3+Yd+vlK182ojrjDRg/LwCu+nrY/0IcVjf+3+XQXWgMakH+b8q5
VaN/37sl+Npb7/c1NN2qE5aXceX3zIRUlwf46JurM6W1FS80+IrxmdT+l6tpLrwK
8Nj3t8FHZaVW0uGe4B5Yk8ALL9tGMH15HfQIioiGiEs8CzbUK1eIsFCO/AzrVVER
GSew+bPMjZrHJDrjXlzAvLeEO/zsbtdM3FyJj7qBYyuMkQqeKoy4epMoNGxtRugD
dS6Q82NEXxgHEtToQG3oLU7Z9WLP6XXaeZZMHw3pRo/YFdKG8fKJKxQn2aUeSxr/
Bjiqqj76uXcTRuYS+TfBL9Rz8fsUKlZtQfy4T3W7bPYrKDoroErkIP0NQ3MGSR5H
leQIsyi89bUQ1JioVDaPotZLA6S32SDu1je2VCggPxJvLAdiwDP8iZPcOHtpQI6C
oEdhNc/cNmaA1Pysm9pFCNvU1CzrhhrQWM5GBZnYF+lnCLw2V+jTMDmL2ol0UGM0
USv77VSb+yS+auPDNFdAT4wquVS/5gBt3xwUW2HqRIkoTXfzkVeInaRUWiru9GMu
WasE4M4AZER+p58FfcVpKKf3B12a6B6v15dZHSPPjbGDkEHXsWRpUeNjZDIA4uQh
qJ+OymFeHRKsoYwUoSynw/wL+yKWrVDZoVtpo0ZXkIlEzfhY/aWwmduResr2p21s
ojTeAiWGm7XBW8U2PiVigMbc+KU7aFOPEggA2imHHaUxkWQgDHT6vsSL8E2xQkAs
3QgYhgiKNGcn06ViSaIO6ehUczOncg9YHuJgX2gCamjkZI3yoNnM0ddxPaKodWIw
sHKUjn2SxTSWe2YyNW+fvsrnoAH5JoMjMnvMVOWk8JBzMMKrikhQtx1GSMDKfAVD
2cZwmUcufgekKv4V8SupBiaxqOy8auM/ke479kMA3LmHKfuZx5Oq0lRbsDuJa2oJ
+WcPAmP1Y3HDUDPVhhjv1/7v74JOvtLWfPwETVlDr7PSVXCVfnEmnQw/g5rKRv0i
D0PKtFzVbfnoteamiLgD+CT3phVgyY1xbu7w90ykvXqanoy1DW4SdHG+/SnIFCFg
NnlFxFQ4sa3yg4AAemb6CKBSaDyIPVSs8k70u3yMGWxOD7xmuYR6OvypZ4a1zVzO
m/V2qqgClJngoTDnAeTHDdTZqMT/pVo+9WbGCz0SKfJkF48jfu9mW2UJQSGe4v5g
rtqISY3G7NkgcNqGHAVrPDe1MzA0ShGrwev3r5YfwSQOAeVGM4u4UoPH6dzXyYBi
X3RuZbgiSm4BCE01WWV4AulJXnV4xGf1aLjKmliCBCo9M0Agc3mxMrCYeX4RCtol
SABS/uKeDlcvBBpIRwrHEMIenymphJPWesPIbVbV/nOvQV/6lS/eKhrVQiCkfeXq
KEH0iah7hpSdTeh8GrMdCaysg6o+YejnrCf+ahf6bdKi/6CMX9cAZrxBhjLwRhqA
cYggpAw7lhrvXmyD0tP1hUUo3s5j2quo3i9i8us0dsBjv8Jr0ckm0uldy4ifjoFq
NEL/3zeejRIA8x6+9mz5AZ0PiaqiPUhjelRM76/SGO7zvJQWAUHfaC/xelJCv0J9
+KnZ1GqQ1QzQ3nqs3URd4ugBaGNeqNBQCCqWA50dscnRlbll1q95l5VId3mKCbhw
lQ+5IpO2WStroQfFgaNAwZiSk019bJRv4d+22g6zi0eEyaYepM7BEfBI3vUd5hv/
UGnjY1StaAbJg8QlvmsOJrlpbnaOcBkT+tbre3CTiUcon6HM0t0sCyZsxfHl2mrW
ULg18HWnfXGIkrM3/jSmAIvFhYjOzBNsTBCPZguVdbRbp0EN+mrcho/Q9Ge65N2S
xyJSsTSDazhUIhemVvqEtQ4XhCnYlD2ItIIt33+HI5iGEpDFrdtVSzfDgmIatkJL
PkXMFoFYBvkIpsAHo5uirlfB3RC24kAhQfruL+kccvATCizHxEt+gXC4aarzPOTO
pFNRfLAYtiGTxlAbYAJA8gm9kw1UaUB580/vZzIe2Mv3NQS0wfQA54pWAEYryxYf
rzFu4lOJsAK000GWPiOAqcjunkq3SjV+NzEbRlLvDaNTHR3yWQzegw5R8+ZXzGFr
Yl0F9PFcetjKzMpftoK4gneeUD6obphg6vF7rdPVCgy/9yKIuMVUXoVOw6D4yHgW
+br1FMmnFgo1ph4qsUSAI9BP1TNwPfwA6YIaWVq1mZxUUaqFTLv89Cx/OSwUTwoq
OVzQ896OWYvynERxqwbGadG0O6Gw9NSllRcOsWEcwMQEcG483Jxov1PxuvNf40P/
/p0udS8ExcqCJWbqq8sfqcciFnOSpaeRKGDB+sjqQ3jBR5DXXIigBXuDzgQDCK2C
btzDc0HobRGUeNDZFVcfXHp6BS7twIq499mpdZHe6HMVnUh6RJ/iU8KFQzRxi3T5
N9sv6T05CqXBz6okZTsT+pii8fk/Qj7ccUJQqSYF/TQGjnmwRTVBVhuejoqp/Tpb
IWXAq51vZJnKX60I0ifu/qK4tHaXHDfjZBbpjWzgbXWJBxBqaHaF+1OUeUVbP1zM
2q8Xpcz5W2Zq8zDf0u0qsu0qjy68x9Dv2xbJrZXiBNmDnZA+m3jTXSiapyQyCmUk
6RbV3rPChGSA2M2K98wHLs1ixCgq250NCsdkB/j7bteiT2HfE2J+aW4k9IYdcRsB
sZoH4p//ymSpAPR5tFM2qWfAh09YHgPYMUu0vUvYu/Rtp552hBqPR8gU+S5KYlYc
evkBgzqeg+jBe0dS1NQ/lFdGYdO3Q2o2CcvvhK594irnvljzw+I46i+4mLEELX61
nXB51jmfZmnhAbp5wyjssBE6ildH5TnUpeIYTNH7seR3JSTHV5BKu+Y072ogoUDj
qrhivQLVEHONW9tc7ocrKSZmL9e+Bt7HW69ZcR73/9CdF/C1Fxz0RJ6CizqOVTOT
wAqoFReoU4ZaZP58+oloHzlCCvde4YlcJcGcmdP67OU3Rem656jiAAEMpSq5Zxhu
ofEG0KjV560dCcPokr2Z+n5HV0/RVD6Lb/aTzJN1SOR8kR07mtN5EJ+PyhlnJtEK
cXO2eUPgFuS+NAlbf/Qb+SBgyVyH24tugMwrizeyGSOS2gQyOoVXDedB+Dcyh5/c
88Qf+AO5SEXFFwhQo5Cf+rOr19kDtxQMAZBEEbG26K+EMkNq+sNzUxcxQPzruEV7
wr9Dje2j9bDIBg2SljX2M28hEW7v0dgjWzwn3k4LjX73H+2BhYtTm7pW8w2Okt3G
d9f+FxlqmzZnhVdyGTwfQDgv4CseCqmeBgb+BOILNhZE8FEdVfQczztstkth8UZi
mcnRMOKyTdT9vPSX7H6CBuf9uf+Cy14WZT41OmaJINS3BuzFCB6NvUoqX0agFKg2
+ErGAyHlNwi0UUZ0hZFI7pLbUPQ6VGa0TD0BpWDYXuHT7cWWq6E0skSDcs7eLh94
+PoVVb0p04fZG45e9FEUaDoBnMeoZ7imSMgj85SglZCYrPntylz0T0OUdzWw/bkr
r8WXTTSaHPG+hUIsB/PNotKSrFfCAA+dhb4n+ymusDymiEFJexI3Vij+FUB+FMEk
DCnOCNb8x9Di8na4fvrYTyEjFMp+XdkPJUyLodgMmlWgtL33ZgoCU4qbv6jovOXz
bKQs4deUb7FGpX5PtDcXFmZGA/1EDdBVXjT+qpc6mgD5dAbemRjeQhqiuFkRk5sv
wSGZIM8SithibJqeffSZ+tB976mB/WBDzP5njVX9vobIe8kI8j/JqwzTWEO4syay
Sy6rXjOy4In3kOvYO4Pd5TiwTNHkF8Oig3TD6JnBzBBZjZynFzs6E7kaKgtR+Gip
2WezObovxgs6K61o7qFU+0HNAfPDe/mXKIHzkx7pyyuCxGxjYwdUpsiI4DywKPK+
lO0+j2B1Ea81FuYiJpEZq72PhC3dJ9/3Xl+2oJX7URukHe0rb4Sld77XdaWa2QeC
NIx8OrPbKBSLBxYi1pJD2PBwpg7TMRLITXkxCffCm/1E2RVJL38KMq0oULSPF5qb
LA2PA+IRd8IL7ebrqlUXm8UV7XkjRshjISYRa0v6n7yqlcTaJSIyWALcu9YVvRlP
bBU+E8/LrvmkctxW4IouQGvxU+8jj5unRfcXzbFGasKR0jXJ0ZXLdWzXsq5/DNZP
EA48KfobF+79a6OOUM+gydV5zDqYTofyxqF4+pbpyQG3BKQuUjz0uDoIQ7JkEMvz
CYQBf7P5qCRd6iPDfyfLs10w1ayVwXAyY3oxEh46GjW8JGWO2ukhs3UxEFV4aWlq
7dmOaQSKrtDsoLd2h2ZOuqxzL/fY5yRTUSGDZml1X8h13oP7c1bosMgR9eO1gjzn
0A8SYqHGFa9kjr81fgqtXlpQfOFf/ehLOHctPuI0YxlQSmETuI4YYQRMSZnlruQh
U1i+gNyWG9RGNWLUaPaQcWPWQ/KFXHGbmH+9tOxYUeJEOTgHar0OCJg2Ryo69eSf
MYehAct4NBBazu7I+popuDoAP7ShU4im/Xlv5LdkL5XtvXUYqN/v9R1eKwX7tVWO
w+DXBL6orc+DtgVMuy7QLVM3kszzgKMu0D9pjxn8Ny9MsrRmvykyDRwC5a3GyIXs
dV9T3acRgwNVcISVAXldBsDf9PNkVwObtTUJEqGtf7rxvoZXgS/gxsDNrK4qnxZP
U+cTfsL66RAFT2YgItKe36hCIYeLg3Jd/O0BTk+6NJVTGk0FfXD6rYUcRJvWgui8
WFRmfIMiDgt6ECAINteGHbPzA5smVzOa9vOVbP8swSzLwkk9LpPzTkdd5QOMKwlg
gNMNU67f0eoz3jojUj+zoKuqoK4d5o3pLdOy6D1BpPD6OV3xSDq45DiFyTAF11ae
4qr66+D1WvCWTTSU/756mvKXBAbH2SdXh6zBNspgeb8j4f7JEFQa42pu1EsdG6X4
9aGj1l/I/ciad4GiVWhIUZecvN3Ibvrr7ACEQma9hHTzux3jbT0MM8RS65tjuJn7
URUUxgd/3/3c+XX0XXY2P5JCocS5OkI6LP4DZq6LLFBPQc0ivTYMZmk06rQ5mzES
9wq+qdm78g5EGhX+1IGzI/q05Nf2V265z0/buQRj+VAd2gEfPibn8a0POO1qtMov
UNB3rU2iNNAp9enMU/PpBpbZhR0kmX4CIfCpEtGhHU9bnQ29U/jKr55BmwLbu9hN
1jxmkYOWHYdLmV2Its+uGkAavwQdDrCALH8hH5vTNam+1IOXch1UHg2qUGbTcfc7
njURePfwiukvaVVc/gYXl7fbDetfKF+YwGrzCCP/n65x41UoPl6zXm8zsC23aiOy
yj3cxfaTnE+i5aSAaGdE9iFOg54EwXAyipXVkAfozAV+Vpp+PH15nI7UQSbqiP7Y
Vi5H1aTALk9C3KCSDHzS4z0JBZnpeBp3wCw+tkUhdy6tT1PaxS0UaVO317gSBmR6
6L18ytqJApl5IE2DjGx8wXNg8u4yU9e95jfXk5kdh9lTiMwKcQMxgNHLBsyuL3o0
yyjSvCoxBdcpCnd2iuuNZC8AaUKT/krJsbn0Q+2NefjhUEsoZPt231hIa3tGhEuV
i3y+BQccYUjPEOeHyXF6uao/aklVvln91FEOdvORj+fKTpFhjcEgTO6IvkDH1gkF
q8OW1KGKNcSf/zgVpKwa6Zpd6VLg2zOen437NP0Gr8LYTRXeY5DX+LvFtyb+zid2
Atz3GruNG21jD4Ux9e4Pgad3LQ0fraYlC7rIzDlDPFCySlsN/G7Ns/xAdNms2dHt
/ZNh3ksiFPYeuzcrIjEcR/nVZzgY5HECvu/7lpu4aIL/gGHkgTcZ0MFp+XilaCRB
aIZrnTpT7yKjGOlPRs1F3RAbv1eKuon7SFag0h669TccYU8WVFobELSXtwQsvGKH
8BNsKdZSqJ8lYHtUa0vstpo1LgsoNeRLuf9AmYkXwA94EFq8po/hs6vA3stJiUDT
MwTCEU9S7qW4+S1x0JE5kHTWlQGTR8RSMj/xCnyyRhBV8Bj24qecFs7PDW3n76no
oksVe2kcoJ9bGc/XUxM7VQx4oWBQQiGlonRiKgM6RpH3KUfLEfGWpKNpoYeUs79/
M5Md/NwajycJ1WUbQEQId781ylR2qs414hzxXS3KyyoKEpBxiad5bjRUxT6KzQ6R
lQuT1gT3TzOIo3yChrKK+C8wUPXw/zBVxvaKSQ5mwheYhxsKIufRz1G055UMzAYt
1OQAwQ0NP3+5Z73XIVCA9SCbXJjo5Dx6WQfLy9tK3GOT99Xs9UJHCfgJEC4T/xxR
Mo0glI/RsE9ew/rp3kBi2RcVqO15yEM0wDYoviuAoo1/ARmQGaAt33A2365qREYQ
gxFrI8+Nuy0VVuQuPJtmLHbJ9E3SX4xsKgYK6Hrn7HmBChnxL81Y+42b1FL6S6lh
WAjE+csmp5Sgbup+7as+IsoozjYBYM/6WD//nfKHx/Q4uV+nH06o3nx+9HacYXzW
H5+q3QaT/U8/RCzz+Pm8yPRwRqrQ7whypSkHydgubFpDlgh0JN5s0t62nfktQbLC
YxLKbw1njnDmRqvUKy7vcgW1XJATxc97ON9JgbUBTkgzxTR1HSNuB6htGfKdTrhe
OyxUh4STkWdrFPCbIHsZTgXisxfLRSkw7qJ90gcAY9txbIgeF4XpumWOrVuE9Rpg
myJd0q/PNK7l1yHme79u72MyoT6Euz8g9F/OGwpSpFvhmHPyL9jKQ6aIRMX0jH9C
nK681T9h73zbSklFjqyGm9TNMb6XQsuCN54gzfSOomYqZvW3Ad2u8CVI0Ca4WLzD
esoN9h+VnWpmnB42gR7DYkeYYpTK0SwQM2O1++eBZgFcht1wzidWVJ1+u+6auNfF
5OVYXIBo87tkzVKltCelnuSnqOzvUMuFEt+zRqdEB+k2UqS6PAa+txMuggyNz4sb
O2AkfNl1oH0yQcbXs0lzRJlygv9IdgHtkweqfWM095/r11DvgSR2FoBEnLiWpG9u
o1/A+XMetWG0b6NDRYKdOLLre7xEzhP1JIAM1W4GCqLCkEeRmXTDgxqvyA//Di1H
dpere3ujMZzBpGlWWf7oLy2FArc8lKmbuM599SmXgj4bL64jxD2IyrcCV69KpseY
w5c08v8j/BJykpkRBosg5smU0KySeWLBo1h+p8hwTmRySOO1YUzbxPCJ8bR2VGWT
/kAljwa8faDE4lmusbpSiYW2WY4kc+4F/kxT+9WwG8B/D/J05kbtHF5AjePsTt71
fPPgYHNcHNKnA8PKIso4zGHXcXyO66zigym1uOotkYSd3MvvPqUEhkHM4UdiMTVo
tGpNqD67zyV7xK4/gDxEWxR4GoiRGZ9N26feAUSrBa6qe6Fq5Je2de3VbN2u6Rqg
ci0hMRg2wyrsQQbbQqQfC9e1xllN6UVfqsEwpgeBBMV26o/GK4M0+Q4cLT+jqmUo
QRUlhdVljk6bSQgEpTuWAHALelXACltuyBGfPbysGufZB0ahEW2LnCmRWiwJchrU
3SPofko3X/noEMl2Koyhbz5tFIHG64b+pV4fztSHrrKWKVliGQNdY5FjCQMx0Gfo
XJrwlLw9agp6KpsZrNhmaRUYNFeBJm0VPX8BdOcreL6zB1Sb6HcEgPyDQiFqSNv5
CUyqlcK3o5kRvePox7fGhpODxvG1zkzKz/UCKIGKhMoHQkH5ZWfYazICfXphbjGS
yNXmRpNnQ0y/RNllY7ODAO9NDzkloci8R3kJAW8s+AEiatT/5UC4JeB0MZEfTXdm
H5kXZ/1d/MJ+18Jnmx9diKb7LLB5jmn3fnHQz8XR76l0QlnfX0dJacr/dpOMhZC3
4FcskXm3FWfKUCD/vpC8fHPf44tkrG3ivcsMuFmRMS5CYDMKy4LcHG8slSYe4hGD
JaO0ESN2MJuMiUToE9i8sG/yCSwKpBwpwCiz4CA3Y+mgi/xj3eCDFRSYmeN5SJ+I
XQvb9FETWLUdV4oJ4bLtT65CStzh0MjyJHzDFliltD9eO5T/NqcIlviX+bQExQ6a
wlqcgpoCVqU7uyU7j2/+C0AoxRNYIPMK60+/b6ueI8c9QI+dtUey4mzPgUKcPTsd
Qkv0045H2+jRF7D2azP8x+81KgkaQIdXR+8rITiem0khmuuRoTlgOX427KN1zeSq
0hrrBI8JJM2iQGajYUvy7YtfK2jJDL88oTa6jL/roHmzbW/z01m/EMW/lhL+nkpB
n0+I8wm3Zwqa7dzKnFnCV71J9W/4tlFryNMqWFZOsIstlbFLDmqSs0PiWjWQqJ8M
1n1IaebZPhRv6Q5mJyQgFGeXWpv8L63u2KgRq8xKyDYFvjFa9dkDp1+/+fwKSHWi
LlIvggIFAdpxCSTq3rPGEufHJ2IHuNNFtqDcRrlS9f4WlCZE1GoA/LHpSO/Jg1IM
2eN9HifUTX8FxXdeKif/8URfvjcZbReS6v3iJbaUNJTN9g50g4piPopTEFhWFhJT
VzY6rcMnikgzvv7PDaI9yHynmgf7twHDpiwqFlQ08kfmbLzOlOJnwiwgy3WVx7bW
FQl74umK+OOpFZWXSrgJ4K00FXCCKR4gS9TR4l9TIxk1LiVNrg8F9LkkY4riWyv/
M+rDvMDR1u8Kj0VsDbbhz9ZdwjPqO+CT58r47FvFA8gPBxgZkUf0b0K3U2ph5nxK
wy8XW137INMZ81zTgHUXS/0rHNzlZC83sXaDKWeFsOD2ZyBUmqfwVC88/gWDZ9j4
2xVPfrPJ0Igw+8TUFbHGY/xduwEZEhUzIIzC8Z6LSV+HHpxMGDOVP0Yyu8K2GjSa
n2K+3I5Bbb//CrZCICxpmZzMdcYGCvF9FQ9IZUSu31dWnLOHvM3qnVrolOYjgud4
q8F9Ys3peGiCbA41LSUZFROzp4k0Oqqm3Ko5XkelnW06fn2E8OlG/WGNttrLQQwY
XK65Lzd20NLjQDvQBw3I9T23BztOqAKnlyah4EnkvbIC8ZEaEw3J+qZdvTALVoke
O5bMEnh+avvF5K6DyZkJIEICmLnriu7tXV+TmtH2qvc7TsFwEVeBf2EileT3ALaX
L3ojp+OLV0iHIBrTqz1UBw+7RFbkJDL3iq9UOTKYIXhpj+xrMDFTm2P3YCyFYcVE
ZmEWCZzQAXD9J2PTuFSZxSkSzcaOmF04H5uR/YUwpVJG1ccs6EAmRPQurPY2wzXl
3ClLTql3+RE7SI6p9dckm/ONLKgc7qPWwl1qZ8jiH7tssewNGwS9T4VF4ySL2vDY
+6Hxx+EGHo2EizHZJZNxNqlA8oCQGepnnwnuyQ7xun1oQh5ARnqsYTRUOBCdnSnP
1V1pU4sjxM1f4xbG7J8A8dFH3AlQr8d8kLhRNIrJBATff0x4kilQczbBwKmdVBsv
KzjsgYN+GzfJ8SKuOEDZsAH49rXbLfSsgk9opojU7VE86pAYqInM0dj1XF6F1KOZ
chQ5e8gWaTti8q+fCxZvgM/0tb1PUaGnbxTCcBNA0WmvLxQvypthuzX1QhHnGRKx
OCBMW5hKsjE+GdUlR5/m253TWuizVPdiNrYdubtycnEii0YZ0KR09AVrctjtT8UA
/EXkK0+EbU+KOygaCvjVXQCfFzNMqHM7RVnnhjYileHHahzy8lOa6d2EnLwv7bRY
U0KEv7e9bC7kCNoASeN0IOhs4NS4VnLjaJdEp2P3CZeq8RsNAI8WVd/Ut493wki6
gBopzF4GZ9zLHahPNH8VYUkfm7dVuYpsgbJhWm0PubWHDSdsO92Ez99mqHty4Yy/
uDOm4bPiIEEvQUz/krGBud9YI8cdmnScDbPhGITKlIi0MSbHefuQ8ekwWJKufS+c
7eUoMSdK8F/XqiRYnGUb/lnyKgs/loGobC6jKn5tHynHCWx7XF5CujXm5muuQKtk
OT1+ovDvFaHYmlyVrYdj/c1g/tF6hud/vqm0IgjCMvAcAtql5A5CwV+5B9QhaNP3
KMizMRCybumwdSc+GYPPOgd15mQv0/jYtET4XliztTMLVPseq/V75wGwdlqfBNZx
dmPFsZeQ06kH1uxmekTEcewX0Uyiw/VJEQcnozACS4rj101oauQvwupj5T3QjMOi
A4nsTH+DZYrjDNlvdjXAvoJt7exegJUUprWi4suvuK/PFtlTth1FWoCcKMp0wNpP
gphbiZ/3dJgvg5hEn4SulkDYMRHq3Vq5Kpz5QyGyUrG4XrYuidy2muV84VHAaMUV
qiQUF5+d5AOKx9A8VjSA7HkAjzN7OB4KGgY0DRJbJchGQn6e10ONfx4jdAIHul0J
flrlkT3nE8qd02fF/XJxmWgFVsPqZaBTrtQY+NSvGIpe1YhdbpIfy3DYewCTlO0s
LEmybkGbzWr8BUHobbNBtMGhlnj3xU5QSD28fmDxJuHVmCEwOw/HOlFjlJ/gj69z
9LMUVgKgGGORk4P3DUagCCe1KYPKWel2Up6rfwPXGAjXOkT/N/S9GfU/9M5lZ1ga
liV24ThLPR8RsPMZY5U7NLhMRSPTouqaYbmMEFxiqVq70LfCtHtIqGjzqr20tyAf
ovc9JGBUz890N/QnpRDmTRXcOXaEwaQ2DxB9TAoDrrlszzJ9PA36fbL06PEpzSdr
AQynI2vRZmjNo2O3ggaHbVSkEadENpEkwtbo4VsBVJfQWdCFp480DwifwMoklwSS
Th3HR268vJgxXiZ26QY09kdw5xb8qBq3mPDB0nqboHNY3qFWniJ8evMQk2elALeK
BTVyf6m4SIz85TVop/fpb7rqYjLFNxsKaouWVDX/nPg0Gn2xUmUbpRB5LeYcZ/ag
QyyL11dl9i+91akfqscaCS15ATznFwK+Zh806Kaiicw0NhklinU8LR8v+X5Ze0SH
rngjNoddM8W8ZmGCecplDrKlP8NRNNk0jRDILF17YiB0vpQg52ecCLZZMiD9zseN
/YgtrPfgYXyu5J3H+i1w3SFsG3YPXwvbeJJfJBT4kTHcfq3zLrZLbdW7axs4dpXd
9go1HryCLiISsiaWK32mwkJHSrwSC2KBhcjLCpKGA0j0lbW/G1CNkBTdUhuD//zg
HpAMCjLKI7PjmY4otdaVa8r97wTjH3HTTdHea4F+8U6yOnnJe6pRcz9dzpK9jzTz
ml9oK9kNu5GN5aSi0ap6Wf5Q9tsysgcW55PgAP40gxYDTpzd/hH5yPeUEN3D1Ppq
Ua3YYaKuIhlnIcChumLrk/bTzdyYPCuWEJ+NYZsX4UDNykiy7cDGfQQdYMhyNQwQ
5ckRccPpUwMMVITaTlZujR56B/N526UGbwUPiHqgJoiSjDa+SmuYXtXyUA+tyBn7
zWJLoDlTRpxo/wcYNmi8UEhVQ3u92K9deo84mEqYNh/OapNtXCF1dOnXDz7MtMvW
xZDdtZdezaHvbnoP9vGBEYO8fN1WTmFlHb86tRRjBI5aXW86wLLirNxT1KMYibr2
/Dc7JAJkd19bCveWwpn6deBIOVHzQAHdrffd5KDEBvqbpEjl1+rq+btXQzJDU2Cf
gineU+ufF/s4OjjO64QwDYzLHG8jT39I2LOv67vbQQnmqrfzTkcjkoWtEKMfEpb1
+hnbJSehIQ8gCIaXEJMm73ZoWd6klmscTBPsiUN2W3KiK8abPxvmzytdjv4GCw0p
BSGpceFB5eu+CjqFfUwAzQN4PmYjoxxLxNX8qJnqPJuUdExSGgetT7Q3OoacQAtn
hqaeti7YRh4iu0YJpWeP76+93Um0Hs2TH5/3UHACBH505Oyu8Qdg725Ot+rHtglx
M6SQGxeGZZa5WklPOu+U6vPViB2RTrv+6ZK+ZGOoJTZ92R+abb834FE2B1vy8CaR
2q4DFNRwiLG1+Ml2jWyGc+Hik0BKHawSAlQSPJb7JSE2dHcD8qDr1y68aN2q2of3
gkcyyQZ9cSR9xWpSjLneX+HkRYLOh6bf0KNHAB0SFoFR5tBj+cN1+jojyoycoS+p
J9N/HHkmUsrBK8QMqKqay5WlCi2oW5cIgfhQ5tC0iCecklNv9syTYzDrhb4mnlkC
xipBIKEOd7pmUksjE1AVL2lBe93KH6+BKR6VZ8hbTSEuFo007Hhhya0rqqDNeily
40bprKcqgNrwW5vMKF6ucimh3HXyHXaHkMeA1feV/36e6EGOIH9dvvyvq8LSPjpX
DapusXnRHpS3IMVzpJE5wvRrOa/mNjQpvMC2YAccGrV++/gOePbW508XkV/p4V9c
vwwc8Ql0uVvzwi9xaf4wS8FX2R4zM+HFhBbkpwAThTjGB5nmp7AKds+n5FxJ5hP3
DtDlou76r7M3iDa5c6F98SGPIm7UV2FAwvjlFDAaCpGeCwJHbT00n3HoxEuw0reD
l/2KEfXyMdWv954U9O+tYAVxr9wilu9apX19G7X8to14EpaR4r0tZbUWw8sL4NNY
0iLLTnUdfBhrUkLGItuRpQj3xAsxtcjOzib2ZHkUKlO6p25sH2GG7Z8EmWQZmNbZ
aMJpozxN9wucf6Iww8moKYBx96y3lbAhjhX7ak349xjglTy3p5FdqtQriImsG7tT
yc3EUn0HaOM4YYw51IHXesLYIJBYO/rXvb8tCEGIiR6X33YkszRJQS7Amvo1xDoD
jYp2BfFl0uWJzl5X0FyaFxPRL6UaL71sKa70vCBKCoaWm7VIF1KwXdL70W8bHFlp
rutdE6pNZQeU+c/v/ptoYfieqkXOLRrMIAO80PXq9VRVkMpQeApSil+gAqja5eX5
RV4DJsXqiWUIONPrkc8lpKpcRG+0YkeC5lKcIl0LtGy2eowN1s8SUs0W7XhktR7Z
icuUkyeuhFd+I+S+7XaCzS9eFPcAWenQpedDA1Jtv9vEWNOEtLWNM+eoC4+99Zfd
fUYjXfyrLuGgfZSD68DwWjQW49I+rJGTh0YWkaVPb8Vs+w4rnbY2+SNXGbXz+MJV
65KCBtalKaL7iPJC50CRzbORmbO9QNFx+oGrUmxjTM1ztH2ukCjo1LxhYgNv4/m1
6uwL29ks+LDT3uQW4wd1+pm5sZD3q5l5xrIvrRdctYMWuvbCJIONShtt4Dep6bLl
hs7Bh4j6QDrG542GLAtag9ISm3aTwtFAl8ZQavNA5b8FxgqCi+9jjFAvlAZU8aja
o7Trodz8j4SmPdTpnV3f2nsl60h4wgtez+Kr0NrKpdQBQu2wlMwF96Rzg3O2ELKp
tcfYYBlxf6hYSvh7vh9KqU+8cMMs+Xb7TfL+57jHSfX7wikcdjetXunN4eBCnRA4
DRYwVwH4L5lNY6UXBZxzRv9pIvpGL+OyZg1hKTiHC2ikS6lPIf9p+vpcM9nZh6bl
mAQeU1qgnC54JU8xirRDBVo7TTInLTzN8guFxY5xTlUKltJpX3LJxLbfLfhYLwYr
lsKEz6x7Ju+TOPtG13BMYQ+lfLD1yNMsgdN6PfIDaGb3y47Y8LHoOYfEGmAnC5yj
RIMC+HvGO89c6+6AtlW5Jbbi1zvPPTW1u70Q/sQyF7+oM3xYW/Dq/agMkO80SCGG
EqCKeKK7IpPTsDW+lTHxNn9MbdknzsHG5jC6m6MyyVIxwiITJWdrJGyaZMmOYsL4
kt7drKgguwko7XvWf4plTjHKimpF4nxEzNRAFepNSybxUwS9vA3z68N5DqefvhsE
kAOfAuQ5MEH/kyEp2s7RXKu9ByXmMBcfPCgScQgk7P+DhnD6gvy7Ch9jzjdQc+ud
o81kiv0PDgbuq1AvuaXTugZsv0DAwpRcNxocA0Jr7yJw6nZ4RUK1jWkaCWf0vD4R
DuWnA6ZPUxEZI07kN1qtouyfCw8IPU+flnnb9ll7CO6VBBFmcPUkFQuVQRdnLUKC
4g3DI1dFxs+020Gc+la5pCIT1RiYdjkzCIqPznYbXlpbBZaArq6vC2Lz7PIP7yAx
eEtV0XLmZhmX53M0ieFB8bC0Q/lEmjtcP0GX1DkA9zDDUFbbwL3taMh7W1kATmyH
qpiC9DKXOXGJ4mUWDGd4Eb9zwJew4qbN9gUkH+Fd3eLkfWiVG9EW8aL2GqZOtHh9
C8q+hEuU3R0+ds4aJRzAXaE160AarBsSgfyDJDJZhKF40NROD4kIwHiMIp9heMYe
FdZOMPxKIS77W8J7IF3iBivKRcQZy1wXEnEQTDXylujMEmHdbKLx65HvYtzQv+7A
MZux/DMxK4hG7HCZfa3cOVSMKlUqtLIesSRjfrB8qEhrYBToS/J91QsbUAOmkHJf
AA8cIUAJd2JEJllb5HDuBPmaY6PTmybnJazm/d8H4qmhWCC8EkLLhYDMEgbX0GO9
dFm8KvQc0Y8saQ/v8qlYZF8xBry8FDrJFIGl0pm7ToBPYLWhqKE01aqvnIOgQmCK
+bPx2rgxhcjGsg/6ryFkrjFwEgo3Qity01lWJ3UMFqJyEnziCyVOOeFswzSgll9x
IaQVkkUkE+aeRPsUPTndUL7zCWxtCO/XW72myoz2mux+2I74rbc6lDnZufkoXyzm
VtEs945HiqI4mjaeQHKGCEpFdz5kVTQphAxT6ZDvDKybj7e3GLHoFH89ZciDVOMc
agGGT9SC/3dC6f8qwRLslst9lPKVUzTiRvL4mHJtDsyW/rrHouUz+Rx71ZSfu/Jw
Xoe1MkYtk0/2b8j+4gKoP/Ol2BbhHNv8z2pz5PCvUk068OrAA/R6wzJsdLUTeETG
2LZ4ygNqhow6OCdHjfP/06vqoSxcsTk8eqyor+00n3ZsTBYZsca3j7ge4hpBAdvq
w0LgGUBc57Mf8MO01I/3hDPht0LMnElkYDIBCemRy6tYyeF0N0G5Rm966PaY2yl4
xa06AGa/6AU6dw1q+bDqLYybTAYlE7GLEuP0aJnCv/0fuue+M6YKs6fii3Dzz7GJ
Tkv+EAargxD9e58a8pY+PW35rSBidazpX3oBidXwDUJxP98tFIbKF4Mc5CbNOnkG
XFYyaAtMeRpiOejZrqPv3PPnlf1fKVtmMlzyT2H1hxfJhg5Vj0xPOfx2wP9Hskyo
duf5XSSeHjb8M0NQh1wgXEw5q6wYk80wDBpETrInpG1IMKdWZwvKkESJobM1QW1s
MTLsiqhxXWQ4F0EPVrLSYkqa8WaKNiDtStaw0xRIUKwsgQNOqw+QCW/AFrYMzUa6
Z72zyAkjWcAUpKAPTMP8xsCx5pudWOva5aroea6N4beDpKHZm8ydSQJNq1eQJTov
Nqgz89fegp6vfMVBtGbysZbltTMoBPy202DBLQXznYSbKSy18sBNnuDOoCIl9Lrm
fB6hYWf+3CfRgLOr2j3TnCocap6/z/CLZBmoSDXe9P4NxU0btbPhqf1efcZfURB+
n70PHZXWuaGz/1hvy0XnlzLx/LxBwbgvdXgScSw3Q0e2Y5aFErU+Kos4aqNW7/Gv
H5JJbgLfSwedqJ0/7D7qYWTqXoQRK4tZmBP0H88OebtKNvjsjY27HQhTnJTUxfPA
CuiUGoavkqtBVCO1xPW2Yys2Faq7rIR5BjjniLngFKs8pUVxZsFDKPUkHOSD3Q+I
ULy3pglum3jXXNR7zG0q+2FVjdi2aLI35A8PfC6/6LwbyVQbHuZFXFYYl+FXMvcK
BykyrAi5tjnFLIQL2hyVMp46Kg07DeFyc3810O3vlRdSeYndtjQUgPL5Q+mtSAc3
o2yBUhcR9lhzxCw+WFj1UPvqvKHdHgGN1wFwJpAIP3vHrMgQuzbUCzS3WdI5hp6K
L1VkTxfk+me3hPot5tCoybzr/ffD71Q/mbXbkr5sVPn/w8eAtM220VKTINPXUhYD
VG+ROJS1hfFBiXYPOacWwtmceja+Z4uwm+3QxrSNL2tmH1WFQaNSR5x1KJ1KOyh3
o6kX2gCZ6+rdfahexOJjr3k220LGiU29sihPkY/V9Ay1f7urw5EVxsU2wpPbkriD
Ukm/nvSazSQGxMiFkKDKja33bQHQS3O1oHOgUAGOdh9yOrogtL7/rVYoc4MpHmaX
gc184o0XVKbrPKxty30franUnkf+gxovts35KYOeWAymS4XNgHHnD9D8AT1leG79
Bn8/aY9d52M7FVpAiI2UtMMWvSjbalboLZ3sN/wfPLPnRbfitBFOxSBBnbO0X/3f
HDyTxReGEdTUdK6kd6jO9htMmdv30Xg/JBPmWAvm3HFtqkLoKluDJciomWkEh4k4
cwfj4gpZ5Wg5UYjaXDUrg6+I+91clfanHF3OGbFFo87dTxjZeIdY+XAdioJrCxmW
uI3TG5g3RiITPiwSceNVJEoXyfx5bEvN3EKfUA3VcyXiIDphgwpDRc/8D1hLMfG1
XbM46XlV3FweskGrBqLtFZ/+aNfkuFH6yn4nP4BO60ZoyJeQhHb+8d83a6kzW1zy
Ox/NA3AzTilbRcyjqsRCO/+zyXnJreUT+w5mo8zChsUfVrZ3rSACGQgnZdMbVPjy
1hKyZkxmy4gfYNKfUS3rLFYFtDOIhgh9QXU30slaaDYmofaBh9uXu3m9B5nuz+V5
d/g2bAOKfGaT+5NzitZAuld3FBjNaSbr6N6/7Zkt0gQfR+qSOmjxRXe94vmED2LX
WbQZWrzbucbBdeoq7EqPBzs/RrIrtjYF5Cu//bWT1X5uD9cOmjuY0jjE0m01wP2G
X01ahxEwUmAg41wH8/OO1lgc2gX07UpIypXVPzj7NfTCrV7AtAbKpivsRuRZ0bJq
L+9M078ddWqgTutfR1SlBTp5Nw54vcag+yXhTf2lbGptI0LEksCbLUCSwt39IIJ6
zQBi9OGevUaPcPsgGEcD6SC/CXm3Ar2byGWC0KRmJNgVpaUSxXg1wrcaUNNmMVPx
kan0a0ETwhbYoy0FmPaZv4y8Sy+jxq9J/omZillOL34CtqGZf6j3/yUMfoVSPhNx
PjmFLfdqKmX46PoA9r7cg0HxYBp+rx7DhwO1s2d+anI9q8X9+cLTQbtFtHiVcI6L
TZHDyZvVdumTZjFe+wpKAPiOI5wBmlWABAgAc3Ui2GV/f7/QxP3wczrcL7n2Jyrp
Wv6fLYZHOufTTLh6vLrIOLGejUGRwKpS7YhVAfXLwu/1Tfb8z4SJa2owzfP1rUHL
dTiaprjtNAQZI2zuI6FSBW1VRWn4xy+KW9rn+Dl9YUxLh68fMRzTa5kapXY7+gB3
6fTncXvb54qxg2NnMXTd6/w4IK3ys+VwiUnRGRVOLreLVAOLtfwWBNS/c32X6pdu
YyUd9ycENluieezJj1oQdTBjwCYUhUdBGmNMLhUnuWCi/VMf3bBtA0+zBLiTrK7t
sa6GSuXFRWRtdgs5w7YA6AcSCdA2dxwHNCRY+TJxkGqaSoW9OT2DSNvNn2YDj5zg
XPCCgXqddMfKgAtMSfhRbVLCD4JPZ/le9XaDxbSwPx5Rrz13IfVIthUipaQuytPh
WkTVnIUQCE+toCj9rHxow4QfYv/8zFFzoLLOPHjobqvwPAWhgnUgGBpaH05AxkOI
3mF+2o0HPlzwkbgQfosFV4otRBa1kPu1xLbNajo9HLMvl+BxcI4c3sLEx1mnaDgi
/F6ae9pzgBMjG8Tt010KgO2zHZkBn3OyI79sx4zToGR5gJmx6yrFOBuo9Ie75RvP
m8Rbu4UyDT24rq/fqZH4LHGs9AilRUK0TvzGzDzUtCWVNo0j4PPxHN6w++weuNgG
sPOuGsMseuFnL0FBgcri6IFB6VvoGWXl1GSc2x+A2eWluUFZTzfkqb1ygMSG4HlU
fL7uSeIH2ic80YLNo/qhBdYfXQ97kogbnyR6S7d95jjkC4CCf7CwBhZKOvDogvIc
qeIa9CedgNlILaHhJ3B9RcYVlYro4BbxFIHXqXwVULuD/b83n7V/aUy+Jw+e0tSV
ohQ0oWGOZx6lwwFdyQ9MBKYQExb4zgFZ+SIWnAdSpXqAst+whgEfoHYZdB0Ub2V6
ZivskcwXdJoNxsn8/+AOwxJRopkLEVbM1rOzCvPjKzcma/6XEA/WN7cmBcY7fNPe
HRggoHP6+i3+6Ioq4KFWGHkYu2T84D3e2jms0nnwophd6maKmhhY7PyO24XRmnQQ
Asy+VyuEHmQ4f+jO61ZQFCO7wur2Y3STPQmmd38aiCxXX1h8cnqtDNAL43Bxpjw6
WRX65LAVa7XMB3c5zxX43Nv6rJBDTOCUP5JpawP3q94/Yt3rsBhpQ7L1BOMieNVq
pLEAWCqrMCYWZ5TMYY2GzKND5WjYdBE3VtpeX5DwZZmg9QshkN4rF+Xg6W+YYNUh
fs/lMJpQ4/weT12LhbKtnWhMm5AVum8Mtnsbm/2xQn7HBWxeJ/A8LHEppPsuleMa
lvidl54g98dgK2hPWharytPPMxMsgI9MDP+cj5rcEp+MFctfsEF+uqZiuTMyZUWR
c7JK/rtO0TZttEcOAxzrn0NHDe88LbyXzr8OHvJNCWDZPQq2IwNrPSFaqHvDqaln
kFDm754MKJPlAdV0IN+tOeCU9er+PKvBmAY5jq39qYaQK5Oz9vM9BZc41xGkMpPC
kRyMZDP+pjkzupStRZWA+WRCkY9Z1WZyg0OB4s5c7VWCHwVXxXcL8SsqLwm2G7K7
2dMenQN9jhG0Pc/7Psad4L8+fOrPWZhEuzHDOnSsLFKc7djn5SAMHwBxUsaKHCtL
EgfujffahNk74nazo/j5kf0zPXKUR0XkEFiXFJ44N3lbm8SdXphVXciZkTgCDtxq
8NgYJo0q8FvoHeE+j53xUwpRXlDL4XwuYbOrqZc1erKlhwWRwcHv+tqm/pI3mKVt
6T5qB6bq/tsqmza0xOi0nWnIpnePP2pF3iX8Cfz9O0sWmDLOJGeOARykoOgn/0ab
5dFMegyHz9ODpwc2WGN6AXIZ5ZrCCR9CSjU5zhUdbVkz10pseF4jLH+cU+LL7eSs
MCy3l2mKTIhgH5eGKroWvhZofIzlfz0bxO34YOv6A/+nH5WKu7e2YvNu4yolAVFm
gMpjVgamXwxhaTE21Nbvzrni7op9y6iCD0XHm+hvNzuefPmdCXOethe1fN1NCXZL
ySHfZehaEbWOruIbg5Et+0UrmHDbWdzJ6ZEKnZX7njjO+C6nPdTDqcNMotZDJ0Fn
r56j2KUYkEJiQCUMpfgcaS1kul8ArJ8xwtbwnTF26dzMGCofVZ4DNruYNXQpmiSi
lXGavXHSPfWvSX/m0GAsPbw1iuNHoobiC3dVtpcRYngxdUTKLqgW6XQ76vs+asbI
ChYEVH+dbn4HKAP6eD/2QRKor0/qdAQ2Gz0lRRns8sBC8OHqKk6MlK/4q4PWgIZY
aG9kzeGDAVF5lCMLPk26j+9wPhBCNJ2edmo2PCtjQPGBSnm7EWWuNZ9pOmhvgrDS
CvA7V2OCLp8BDxnciUPNFNa+xDZX8o/tuvaeccnL3B7tLmLNyo+vBOYBemjQ9PRP
pO0yMNuY8huWXCK887iN9H9POMdCIGeiNvvqzy43VL6lKgfmMTXy0SyJ5QVNW4+Q
39NRn5MXL4KxDLmMw960vNvF0fmb28U1isIaqF56X1FD0w1i0GVjVr48WmzPlE10
pz/awxYM3YzlXaas29+jcmdJkqZDC7Q8wj0p3AWeZmE9LXu3SE/zr3XUZWvBESfe
0ttYyvj6mvfq5qjY7L0y1pHwP+sfNOg/9y03YMbj3VDPgrRgzcd+5cSZ87fVe57A
XZTyVvvde4pm4lnE5r9n8QfL/Gm02rTID9qPABjpyDkaXw+RcU3pvKWqtQ91SuVP
FHP/zQfEbjtLRXjGJ1pZz5TofgvIHvzKrPMDxBZYYuE/+V0R1rfExNMb+LODpdAL
1xnL7dcvqAad9FQ/v5fYg/W9Ecu7ETE7wupJcXtSqmV3zE+N64GcYfKWDtIHdtmJ
TQ3D86eh8TcLgjqsGV3lZWZiLd9J8WsJxPhguuMuNRmLsSlt/cXIE/sUSUhAoOlQ
0I4pTMNjgoN3cRL4ojtFU+q4yX1TUFTKo+qlQYk/rN0JO+WPRAlQ6UBdlHUayR8A
8MJqPwxWEIgD1lRh1Mjj0S8xdxFsME9TRdB78ew7JCgq0Qa9t3O5PUuiedYt7Lyy
Y9KoPgkfR3ieW2ERWicGbT4/tKauGhJQB2LKiTcw9l35YHdtuHkyan3YVIkC9E7/
brNWo4oGNsaC7O3THWvcA1Ge/M1GTWljgtW72T5j/587JWV+M4v5EssiyEQx0kfs
nTqX8QBU0kZYHSYHvz8KSat4fly3ESDrne9sOIf20vx5DuE032FOvpjSD70oECaq
tl4S/lbv7mLO8a7Y38rSENDgBAGdICvVEPc61zzFkt4G+F9PrJRoCl9jxWgtlQnH
Iqi3j6eGejQ9FFDVz3LH83rzc/C7k3kbtpO121cCtU8UC/ObOiF7bLg/cawS0yHi
z3txEKjUDPA5SeucpWc7KvwTtf1PTFfVaRqQwSYX1AEIcLThSXFXI6eNVzqCxxND
6hLpVqRPIkD24v88Bp0SbLLlOHpnXTSbgclyTnBQ+e1McU91JgnsCGUm1npBNdcp
p8ARL4Rbau36d9jgxQ97Q0faK9OtmtbWz7rfadIIxlX15LR8npdYsCQFIBwx28h1
uX3Fgl+pEIwE9VvdP0FuYvy/fH+1KQ2xH63C3S4Cw0n+0rymmx8OY8sVNdnSgZS6
mh6KLvqdOe1uT9/Bw//CYFBRbGZ/f5FhGMB1wlJXlLykwSn9E5A+n6KBlZj1rmCz
0KwL7P3anGa2FHzDxZQhJ+GrUmEhNbak9ql4RMpwl+n5Vfc8m085fPBL2LTNnTiK
vL9yme/0T1RR3f3E+jqROV9LbCIGG4Iuc5+auzDtvVOmPQHuYWCHs3TpTR+43wK/
2P8Kj44G60NUGk3sIouPvhTAof9QXlQ770pBTPvZRWb8i2YKshLej9mSptPotH7Y
klRLpoXIxk9sLUYrokWn4/PwB0rSoqLV8Efqz8oquwqOqLiL5DyKClKrUyNy1isS
5MMDU4GI4qmjKd8V5iMTMwKKcQvr1kPydTciQuLN5/zennKQiClXCe3pEFc37AHD
WFZ7/lAgzv46/Am/Oq7v7xhaYVzr38pzjzwb97glPgR+XVzhS6u51kVugj30yxJM
zEWxu/gRSst5QPCBzc/z4y5fdAs6TcEj0o7VMn3IX1XOA05f0ED0guKVLjd9j/gH
a4kldB7tqxEiRB1ZZYtkFlKP9v+7pEREtHiefiSxwhYbJ+yn7na+QKDBvaC95CcF
rnyrEMweg3m6p6IvS34OhamEuzYDtQLQwNwyPHsz8WL5M3WEhsmKPKX7YlIF2EYG
hXMuTSta3SH8Jr8rjfjVVRQHnBZXl7QnaMFgke6TUdhNsrl4ko8cXOX5zeR833NY
wnEsowytdzsorCYuUXJQhMM29jOsVguy54tgS4+BwJDyqpZbmlIUvO4ieimY9iQb
TcUcMQHCn/2Qj3JR0gX0Jqwm3TpKaYwzMBFFH5yYbg4uP/F8tZQlgPqftM2YYsKj
o5SMjqq97rv/PqoRokoycmwYCy87na7LztauA7HaO12b5kFJq7CLdTD3Mb68Ynn/
0EOAtDvor6WLJzezXyhiendwpdiCfP+UK9wFSdITFX7nIh/wg+07R8hS2ZjkY24k
qAgFp3hFMpvBEulDfmjEOPOLWLPN/1e+oD4qPCDHY8yT8tQ6h2NP/U8gKq+rtRN2
CQ0SffBLHjkUCsQz0t4HZbpYIPK6xmGlJWE+P4fc69Axk8RNctn+FJItK+w3+QTg
ekOP1lkv9GZyNxas1g1fW0nxl3Or+npNWTjxrOYjkAoorfnP4kxIUSsOcJWkvfyU
Qihub2vAe2UJB52Q6jwt5C357/1enYldApuMjrisnmefQ1joBXUN/PtZ90j+P+zK
XM6tjgsV5Er8p6xcjUEzK9QGwjh86rPjTf15wepq+O/5/+JMVVDjXnyy0tdd0moB
ByJF8i8hxV/dK9n1hVb2kd9im6W5QucZ1gEv7eXZUBaQ08kVroWrWUm1fBOe0YJi
7eLJHBEN2fF8QidFWxnCp6ojn5BnFbuENaS9ETuVsl4QZaMIK+GnbApnMt+cYZk9
9BGBqJ93W9gsf7QJswwbzDysCl8mXG/3Suuf2auep8EkmZMB5ZY4J7uwk8zAgcex
Vuo0zS6gL1QlZg/CL0orSqr2zwhQmfPKDF0pm+FPBb3/xxMSZhDzdFkVA8wIf8pF
K1UwG4Jbh6QqSZa73OKxEMV6S8IDDiZltH5binGEwgYB/16aPna9e93GJI/14bkm
WWCw3arDU+52mrNmZH45QrjBL86yIoHLDiAqUZmeuDaoTCIGFy8HB9Qe35RE0jOS
NSgGTyklYNxocre9R9rtBD3R1a4VduWKA314DqO7NIEZ8g/XjcR/i503lgFc20T2
d1SI/i3FoNDaSwSsdh9mSt3DD7HU/i40NUAq1eJhFFnzUQXvltx12J40jL0MN8eW
5OZOUxs/rrVC+LVGv73sPq/CXSyLnMYyOorYYcCwlH1dX11CEAq+/K7oliPLT3JR
slyQvCy8bLqpX2ciDwNb3BW8VvPdcBQwrq+vLKspl1Mc3d57iOHqrLUKMJhpTLfF
8IPGMo4YaUpU0uv1vT0WbB/jss3cKnT+rCBZWdHru6tO/4cVC+FE31OUqNgWFUsa
MUkoV8dD+9HPylC8/MpFfJXvbv5yI2mA7nnCqdDfhjXen/79LdC3cFDCaK1yg4Sf
cQsWeop+BinAdpu9oNLw3vqVaie3DXlCSE0PbxLcq254rQGhIdZ+AThZRVT4uA4g
MDZt4BiHU9g0tY4Vn0vJV7I89Uqj3xwdDMQnFbbIqi+21onQpo1VwcET8B7/umEE
LtkbeHWvhI/LQ2onY4aNBZb13EXhvpwsz4C3asmcYGT/BsvrvKVJ4e6QKzCsH6nY
zi1pEv/LG1uCbY0QJJugGOIVMuasHG8VmdQAvcR9bm/2XPbbNiHwlq1h1fjHzR89
laWZFkADBk634KZkmWwBUI6K5UFdoaq+pFVM2B5E6UY/X3UK1w8mH3HiwiuGpZd3
K/mb20X5xl+vsJbJ5RTwF8V0+afd2XAK9/3YOG5NAJTkQ/apRkvx58UFJOyT3TiY
IiYbiQR4ZX2bebskVCA6Yxmc/T6f3+jWoxjwj82PVMQ8PoMNZU/9/X67zzYblH0k
9DbSnO4PnTn/FMMYgG2mz2UPWdNw9qvqApc1Q9+ys5CAvzsqiCk4zmgGkjPUZI6S
7nkmhE23dwZmTV9XG2iI+RIxub5TPxDYQrOmkLc/ym0WqzPTe73bAhJlE1hKjVvX
IGzNR9Kaz0ZOQe7K/0TtG2Vh3imkwfzUScmhE6IwrmpFvsYNi6M2F2z/F4z0hFZR
8HG8BvJFccPKRi+1gNIzNJahXsXc4mjz3rbpsoP4W3Yr2g7Hvo+iFucyq17Yo8mp
+7Y5neUh9BxULb3+Y5JcudizX0Gr4hsA1xqgi4iU2IEpCoN6uYQXE+BP6o37dceH
3PV8Hy5Isj5VzuxLGTv/1gwQ3SpZ7M3iURrwle8oZDbN1Q8eu4VPHn4PcZ7aWWfr
UPkVeEXKakq2ori5ZfWxXPkdpSCdJ94dV6S9JZmiyEVKEFDPwysUxICxdTNo+PYK
6MRFTYWSY8FQjm+DoYNt7c9eoLU7u6mAg8PgZJKGHgZrasJhwwdAevImGTJVq+8t
vTnjZImDvuAtO7xlZV07kvM0QmR+n2LBi6PMCvT7dcBG4I7ZSGaVZkTTbyABoun7
xJcs8ulVZEuodzAm28oL/qqjqXuiphyPUOS/9qVj/J86iWjZqML9tYhy3J3l782U
KXrtGfzXianusuUShkEazh1k2bV7YTjL3+R4oDekVN3krJ2vrlB+TilDeQc/Ot3m
OL6lNAVD6pdjDnDnE5p/qnMCGiyjnjQzSVy02e/Pt5IdamzZ8i+I874zfjW6UkB5
8ropX+TMaT1u0/Nie5ZhOJ96G0YS1Zwr2L6MAJurkYznt6Z4eZsa6H1c5d1T35gI
+9DvJf8bBKGa+QyR7kXjvG5c4AeCsi0/9ZOJ3hPfiFGQ2J65zRJDAw60rQmsOL0T
WQcb7ESCqAF9dPzEsQlNwEX9x2rXHOhDgu0ak0ukd77RGvvHlvuNTBp+krP5YUfU
+2xZtY52K1sIPtAJsJ+ojMKYlsKZQHOswHHvRUJBOldM4c4eVQbk69X4TMG2Ye1Q
sU1LgJENltiVpPB9SdtdK+KNxrxVwWS/jFbN7bl5npPypldBBI6wCeGBMTKeE8rc
ccz8WoWReQlfId7Rw2UODF5w6Xl8HH+MrHsLTdhAa4BmopwQ033mN0gmybyRS70l
sY9wicIlPpu2BgORw9zFIeyK1mrhefSOpeJM4HIdx22jDteQ20uoj+wK39v6n0Cq
I2Y3RiqN2Nx9KD+NfPIiW6mbsrfCZQPoQJR4GhctQBB+u7ECMAdxwDUNAiKEL2LL
DLhoLNm3Jw/R09wtifC3ZvVAaJMM3ICYVpH6odo3ljd5A/ZV+OChmUlpuX1i2Zbz
XIOakjuZCF1mk6DZthX/BfieCa66f4GjqYXAhPB63n7aQEytEiRIn0ZhtEiYWlOK
F5uuuTPgNVzS5Zqm4lCnnu7Hhu6U+iLzIzAOJ+c2ZAebqESLS+gYZsmYCLORBm/w
GUO/Jaz8ld+yIqjVqQGEwIwb4qeuJkeB89/a1fMF3ylmA6uY3IwEZ0acPsmicND2
ZIOTEwklSyL762R/IzkWjxWrV37eUIqUS7gfE2iG8YVv+gOE6GKbjnO2cUWG3uKk
UFiI7SVIWrrZxLgZvEUQuS+rXzQUmHbS3DBxz2n5ntGWQJXQUW1GBnv9/kmU6mHy
e6bjhfwMlDemy0P5FQAbhYOP+ZFC7EBjWHpRqDOJwp+zERQK+JtFWmAIoxbuG1tH
2OjtGV3S0xHbWO1N1mDrq/fbQpvj3OByWO/6He2a43KFwMZ0uLoBj7etaLUXis8N
HC3Hd0SPpuhQhbOIoPPuaWyi/cFYydaGXOT10lIDIRYPm4pLZQmxDHcvuvVj7olm
jQE+DTEuk2eZfg6fLXEwDVj77+JVWr/86YRoTqPaw7WL2R65lanqGb1OhyWWDKvL
5y7whJm1SmbiHVHkoojkDEik3OpkQCg9ENieMl7qagSrMmvLy/XvcZJHx0jzciys
J335b0MGvzvtlhQrYXqCUrlqW2VnZmDO+JGxGA6QrbKZU4Ec4wL6ePMLgjKvL25d
xBBmnWgw3wSKtNWFQfP1wl9/rkEvTxoapW594m+YrEE5Ll8rCxYvTmNdtxbsSy/S
z9e3SzrA53TbUn1JRvczzALNmyRmYsl3pn98Kvkq1qmQwgqeoMfx+3VGE9MqJ2f0
33kXU/22taf42FnOoCdX6JloiD8Yd+tp+fzfA0V4kECSy67Z+oHF48p8MS6hwIov
BQuTJtI+eLBK0oO+4zZ3pm8seVUuc77BJSVZLk/OcOrfVq6vvhMXWDkUWOw53Y11
3Y0IEnJj1hn7C3b2c/0jNviR1L63Tg+JXlq1ze+GtUIb6OlJWr4vjlYgI2L8kLMj
W1AXfmWI8c/4nd/31apWWCySk//s3ERIEfYUNexnIlxpDg7VRvMowa7j3erYPV6f
0ktUFxJ8VfZHIjfRcmLlevfuZ9Ux0XdVWER8Ygi6tko9koMUcuwF+esB3/3TQu00
uAP4FaJEMzVESWwGiBBxkjcek+XIO3msZSFtI20xAorL33P8FRWNfbEjX/+Cvgwi
pLP7/rtsrs+j+K5iq4a7ZQwxjmB1ehxpDMZj5S1sid99MheCfU0xL97nIMTYckn5
81xYuc7V4HQcEokrvW3cQFdSAk3rEIydCBdolfwP3nWa0OmbwGu/ZipCeRH7HsUv
aY/OJtq8s2dmIy2wbbiDXax2usbrshUOJHXzfKeDKV1gwI5SgxbuvSIGZOmTGT3B
5fIwhDmWKOaMOwXv/jvUoF+yate4UGyvwUI0zBORYjVOtQjwhTj3ZrOVH1ziyTqQ
pWr7JksWjYZJjYTjYdyXEuiah1B7ohCpRAsH9xm6UQtBzGXwH949v2Pcjfk4z7Mw
tz3koDZMmY5cuTrxYdySclLOgACtmvsW9axpQNDNXFKcaLp5FR+Vw2cMtHsoq7Eq
Ylo0/KA7TIIrTuTt/PLgH6FbS55+S7Qhrl3UuoVTPf/tpS82SypYUhhKhqIrq7Bo
nc2LLD8d978SBul/adL1/Ldud1Ay27xx31U0LEnB4jtMBNjBH69JHR5iTMrw5dYx
3KbT7VBXFWDiktitPO6B/7SW47T/Q0cVHffJEU2pUYqjZIhQGXHVZfIHRZ2h0gHk
A9be8zFi1xhgImtDYulrMuNZsnKk7iqrAkgFCjETzaq7sVYwIW9nAVBW1LzqRtm2
xhmBiaJX0yYSHbPKHMJIjZlLxIr1iSXNVR+pKUDqJ4Ibzvo5V4q/fT0wFVEYLfiw
ZvsooVZ3Oi0P3bz04m9u/gh7Zvpq91h8udRSWUMPnF1dQinCouVOJmXIHSw/MH3y
OhQZwyOI+Ro8bXCw7hllYfnphgENjiNde9ESIseLXXKzOxMOqrJoegvjL8vvfjtG
Qeffzoxw4RP3DWHRvRpTowhAu1xaPJzKQr7tkKUPGyMZG6bbdGSYKYKloRU/KnH6
HQSDJZt06t4OsE2fiTGTxW2n5rFwcVQSy/EQkgNbmBjS/jc+7fIZtE7ECDAbvNQk
aQ9hjWoO4hOpeRNNnYT6Eqi1aq+FiRQxqVle51GAMM71fqERScm+ueZXcApUwtKE
tEhfk98rt50amaRUAsM2lt3GMK52OS/sBTVVMigKsMkfHJB665+zwahJHvsMiGY9
L3fBAlTqpwdrQeRTHOOLqWEs94PZTlKfin/2AqPm8uMhFa/sASy/HMrftqXIxC3f
h2hiZXT5tHjsBsrVA5q/85Ne26aHA6YFKCeph/zM2Hb87DxKZKX1oE5PBh01Q+Nf
bvVGrm56CX0QHpiwIUWzKlgQVT+Ual1s0Qih25lTL/TdddSB3Dx45pBaFfzmvmAC
f7NDCZ4o97C2TEgPnX97MO99fkJsr5I6GrHAvKGCLXlegAN7j7nMHbGyTxCZImUe
egURQwUBqo88uOzoPTUpt6qT+HxPuMbIHvzU74Jz5c3uj7ZTEUZdZIthf8+FbAUs
nqerRMT7+1Fq0na6Awtbae80vCZeJNxa3I/5JS/aOjnl6mplF1LWMo8pjoKDASdf
eP6MON1thWqZGVuCxhei9LLCEh6iKRYfp3kZb2pOado3TuQ0w71/StoMj1f+lzCE
RAV9AkqE0gH59eo+fGlBPEzFGZNt91p+0d4vhk0LBFEI5JEs3rXoE6md7KxBFeK2
YJv9MGsGdyYiD3YJaj/hQ8qT0JsabGgCGkEhVv7R7mSyaPvlw2iNQQkfHi/iK826
BgklOIduPqiTH9WoSLCpHqO00ABCX1+MjOEhkmS6rEwilpYONHObE8dpXLcpEHyC
PzCa//GbTNVEwvvnT5+tIBblPKg9SkVkg9tlQyd9BkskMq+T7Kp7bSntm2UHNRes
2ELAu2JnxVC7oDrttCKsH1baG3zA3gVChPYvjKf2hmO3FxF1O+z49+yzg6gzHcwT
8Z64Zsei4OO+k7uF5gavv6n2JgRf72vaLSmf0WNySBDfBvAntmBb2Mvy/xrZbJcQ
Pg7QWTKifw1TaTuKOpshzRfwxOtm8fruqiI+ancpFykHvGT6SWaumBqya/qn1ywP
5EX6XoXZ0EgX47LsrHyIiZtNaXsrC/7ZRmDyJg5PGXkImVMdkagEoUvU8U+K2PKb
o9Q8y7S24RgpyuO5az2ZC1g2KS2RbGLzB4/gxAyjE24olaqA4IC8KR5GNyI+rWiQ
8oU3XvmQbTQgd6KRojNCwoU0txGfe4AIaOayst45746g6Xh6n3RExc3Wtu/0fVr1
qU/MhB5pqCmTIcop+J20ifoZvCCUkysg8L8/+T2NlWB7tUbm731wbe91Bfh4mMgH
iTroqC9jD09g9Q11l339SGAjdrFGI2GzKURwwB7YjbLuHuc6WtsvbzsSWihXjdNe
uErCyF2ygBA9VAy6j1t8lStGV3asbGuii8YDOvZyuAdLgryMQlI3boQKrcUfuQ6/
MTSSTCkGh1sJKe5XgIR9uDbCJEiG5sZgYhlAFdK8U6DnDDlEWkRb8H528GYSiHfY
CD3hftFB7jcKybQyNiWLGA+U9gR/Txjp9aUqSRs56B8ebvR7IbGpJWs/Jdt8WHXa
/dCHgcoQ2Goe8owPAUB614x+lmeGBhSV3x/Bi1X31SIovRUCqlTt/CK0naYPPoE0
Fjwhza1VEWxrd9dwUZfm+IVY1hPP9YDw/n2Dk9rRfiNy/h5NFWCtNPPCBE6heAe6
yoFvRBCJHDdJEdOBJAzCxh74Xnhe3FuIvzatlM1fEIYwi6U7lV8PhDLdGoTEISxQ
Q5ytCfaKEOObsP0HoNhlp+Oj4JWg+GHUneKKZb5C/UScsdG0Qu72OugGflEx7q+I
leb7r0QtOJ/602oBxn7MhGi+VzaXSQpxl63AHtXQz+4TcJN83vYwFkv1hPiHwOEr
ftbKI40LmcQW4b8sjedce3+8tA2OJysiGSCthTtGXF9iGcuWnGE1NCcwJ6ygN/Kr
+pu9nhU83Ay4FCCIZsganzVn7k49kIbR69TCniwlz8XwOT2ezybmDoZQCOrFRQdQ
V1igbO4kZE36v04z1fVWyYAyn1kbuFTRnycJghZbjJyf3h8QxB/+eRl76dCoOo4s
UiAY1se0wU8YUXwJ2xer7L8qc7lDIx6disHy4GkB9MGQhywGBgcj28/sNNCts7bl
pKYf4of7P59BOJicz/t4C8HEZ6A62TfW7u1reE5bfEuxMOwaZV47RLZPtv8eUfmz
KMAkam2iQhEiQpUE+4m0Y7VoYlnI3Wfe+iyvdCX539+ctRTaEW8/C7TeW/sa5tXV
Cij9vt088DS+ckyCnd8hL+clDbejDiUxa/9qbcyr1zsul8AZucXu4xKh2cf1NiKt
3UvnxepsS8QeQti7wRpvrLSKKqRqvPDMrdCyn7qbiIsYbhzBpU4K9VhiZesgoDJf
BN1K5lKk4sdkNgDksXH7MAQWn9LxJuQ3suPxgZWhCtleZvZx5SIomz7+5ttaLy6K
zo9BzaO14goCjpxm2ctEQF9zwHNgD9GlJHCGRFL6NEVDSRCAh/TdI9INQDRDHoz6
3r/Q6H+OkZa+c87Jpw14ZaCCvCWZV0GyIEe3Sk2KUKSmIY6/OHvSriRvEKn9O+ba
kWq87G55ftbFXNKjPrxBXcC3vgVShikocUB3B+k71mJyPQkQyCpGEOotC90U3RFX
5RfelgSQ8G0JCDYmYcT127p/V4jdi8jyp3ScczUACw8D21YSU4sPww6NsjIAPFbC
GVi4M8Fq/JqCNwbB/DQH4sd2FwQtvvboKGkREWyzn96cyoJv8+56Uq6YVOpl8UyZ
DU48bjVv4qXSyiYPYcNnIY9LXZgnNJw3i/D78bGd1VSlO+yPc4DgtmRF/cJ+9cnE
I8pIva6uL5RmUHUrv+yvlZlSarZi6Sr3o8K8b9SrjFRAQh2pB6jgdCWC5UOEInjb
vDIDRNBAxz89O1Zyxm16KlYSG0Ru89wBEOz1kSvMo3T2fchsxduFVtJke+z7LRgd
ig3mh7J7hOp1JFDaLrwnW/zKJJHXeG4c4kUXQyvToiPL7uxclnlB1eq2NpFL2fee
nX+m++P9UEycyp6tmKiaT3NGriv1KbwgtFUI+7DKQl2NTGh4tu0e9ChY0+pIX6nM
Yd6BWLD0PNbGkrHVPau2ECSSnZKcBJC7WRadF8yNdqBN8+Cl+Ih9mjfOoiu9EGA9
3FaVGmMbBdgx1rOHxN8t5Q7NIGZtadc/RpPT5PwXOmxXnrf2TOfQFAyH7+Qu01+c
4s5KRvIcPM6VPmWPZMYZbpDmkwqA0qVj4CAzMQ1jlmpM/0x9QSQawIQDRXN0p6Qp
N6Oon0U6HbrcqP2Wq2ln51e45Ar1cCmHPJ16gL+iMudnWOesf39mhisiEz1Sx/F7
iSnCqkAsgV48r5a7kT56polwyzXSuV50kQ3fWkmK9EFx/fCZ6CKO61QBajh/6TzK
QEweyHHHjJiY3yGsrg/Z1Ur0DtSlSbaKZDYT+C1+rbUtmP5dgyC2uy1j2N49PqIM
R34pvdrZ7jH2T1KidaXje9ub7E8psQU1F8VqWKdM2G9ThteLyfFe3yloEApRCc7x
Lh9MJvzcDaRSU6cxydmmcolz8+8WDcQ1D5XuX/LZUMc7GcyYAJsHZ7uyguCNS0eW
BvmKApdLD53w33Z4FJLh4MnD1usQ3ut6oR3xgsxLN3MStMF22UHExgIMhkvXo7zS
w1jwlFY/sMfHsZFbOvOGa44ofcYJFtxH45r2BrhyZqT4X513+HeFBP/fwoEIeD47
acFiJVJmdnYN5sxMcZx441sv7mxnYm3Tf+Z5FxuB36sx4GsAua94X8ihxrl4d3VX
niDLn8gkkxoG2psKY5oDc5hEhyY09PtrTLQTae8mAbE4lHWEVZmrRLo+55mK+xQA
V4z0c++OglbuPDRB/YYZbNctAic6ZrSpZy1ZwlghVq5I7XzlTEnJWK7+uP4EL+eA
xPDFRQzYtDQ04vBdZQjxFHmatqXr2D0A+oSXOlMomftyuML4uUJ/vvEwPP/ecXEK
0VmGkPUoy7l2yn/tH0D84tgQDxua4J7oLVDOhLeXAzsKkEyTOon8egX+J0Lc4D+t
c2OB+Pq7MopU9DKuUDpnjFFWYlck6XGKTTjny7+ZMsH+0mez95XAm5rGTqYpCJfH
ngWgfAEOYLtDKN9oqInM/lNK5y85485DlUyu6rkwkIDdrWfVd5DGh3RLPMaYeeRS
WRTRaTwtQNfbb5C1TnFCBy0T3TZOdsbZDzitiLBpT2bHDqifvcG9/WOaBdAAYNrO
HN+awQiOoZ8HKgC6nBadYokeVnvjfoCoggtvWpkbz1J/56KjXbBDpi9reIuXoV8G
uQ+8TBBfTip7fnVBQuwFiODTmEHeRqWPZ97QAqRPs7vFUt1Oqww0az9Ub1lskNi1
OvnydNMhETQaHpBwDZxevO5mC8R0DkS0jiNpMlSb7mkEWZgSk4f1nLcLAqGofj/e
cICMFQ2KrG+nssJLs833IqIcT/3ovwvQ+4uI5OfTEn0f1RID8MZk1ah8SKEnGofL
egGVWBEjBHL0aA19qjb+jKMyPX+cRf5q6iAboyQzChEiT9hHxeir3ZVFC99eXNtb
CmMWM9Ck2WCwz+Qf61eOIv/qzBPdbkQER26ThaguD151HM5FkDayQWLtFeywBsp1
HfrhlMyLgmL9wQTTNSMN5AKZk1k+k9LexI9mumK+WiloXO3LNZTX6fE3ByoPkx1h
ZKG6HJOn8s9fwXGmrlAjg10Q7BlgZryYm7Vn7JEsNvb+PATvQCSionWwuNE+5Oko
kpQNV7bntyaMPL8g2TfYR92dniiCqXW5EBe4olOwQVojDffM+sC3yU/ui640tKAe
ID31XW8ghkP5PUPV76NLXjPFOS4NCd6jDwrB0LTN0mr96lqTCdegzGqy2rGCAwXx
HviPCwbGweufRVIjAFqK26VMz7EfIiPMM2LojF1BxQ+7EABO2QDtwMnraFT8mFPB
/uhH+1wykiJFWV1gJVkyEZH0DeCJ2RM5EioYgecOxISN+iQMhxfKavfCyoVd1/I6
HXR/zQiQKFMIPD82wOKmZN6R2j7JjTrbayZiWAThnj92YVBVR63BUUJAdnZsm0lI
A5guqktkTm9bLtKvylCm63JQolZ2vBfUEUIiFPI57bumbewblNzijSs8tGBrwkzw
njsf/bUjxMX4v/aDYjMOcLQnYIIjLbhYhDwEeE+igoXhoudYOn7qUlLdjPhhaqZ9
oqqYB75TM8FLG5vLKok/cLtPlOYPAMJf8GWa1n2DD+uehW0SWrk4vb3iI9A0PGMV
hcYdDlOsC07k3LgKY0jyfe2eTt+yJclmivGP5V6CLAgIDYodYd+bESjr7O7iKcWg
inXFuW4sdyTNBhYOwUVcJYzb4gJvtDGpdC3Z1u9GyyM+ywQisV9QtTUomGSy5f0w
h14KPnWxcNn76cn35gcFoZZVZ8J/8P19xsyU+rI/x0o5og27UiqFGCNaYxpzLKUY
R08Q6yw/R5RooJT50+oIEriVJeFaBadt4pnQ8VYQHObL6PtldFGt6q06PRj3C/x0
n3YCaEWScSEduw8TybY3UHYZ3Gh0euxC06Z9AZBPQfOIr1Sq4UgtwnKYOud1FXyJ
lu1P+uqghLalSvn6s/Nvd+Eedx7P83gZvKQ3cEeKo0EeWQrXiaaCxI5a0r1tBM99
+TBnPaiKs4bTu3Nt3CTc3iSprjvuJwa2HU4Dpmbgd/ZYO972NRSlYqBV7mq+vNWk
+5irjevn24psJbuglJXiIz9K/q1n1EItHGOYK0NpHb9w9As3RxaIniPQRco42tuJ
THIvjINjoYWeQ9dWFYj7KOgHoVymQnGQ9LtUGvARu0LQCJzN+FXBAjzTPEceZkpj
kdSKPAiR0u0phY2/k6HWrTu+i6nod15OPNnz+UMcXRKujFJWkokGEF7NKQf7WO6c
EIzHVrh8Xhd/EVLnkKqNz0gziiqIhiwSxTd5IjAE650Q+0j4rVSzHXJ4aod1TtpZ
67rFZdvQAxzClIdL8VoZNEyGPtysrMZHrUUvMx5mPvn0gwHMJlDhGDWB8I3mefSo
N7xgCq8tMej//HXJ9E4racl4xbEFGZcwtcJ7zUw1xa+O5Kam6Uzv0pz7r1RvkmVi
uCTEgPrRlMt0t7NLqwbMmkGp0+j1Y3gbH9DV0u+33/f9c997yM6dsXXpsUAr0XcB
W81gNiZ+eyC5s77Pvc/NUtOLtgoJHrq+lwan9OjyuRy8wm2z8WZewt4l8d9xrpAf
E32btO8/Q2qjBjrKSlyrYq8Of33EawLSg09l32mXkrIVxdSjf811U1fdHP08Pkyk
wzc9PxOUFepKgNQ1tWtH8cphRHEo0sZ3yHupfdJIXyjFSjKShcX3UI/2VUpjwcod
ZcQliz+iqKWcas+5ZRg7VjSLN+N/lbOMefrL3apdcM4TuefhmXnes7/zcQ+Gzxfc
KcXToIacnKejD3nCbueGIomLeKa1RtYoG1yh52kkOYD+G3/sgRb6AgIzYU10fuyu
nVP50AfD/3SsachIRLegtcimn0JZDKA8ksQq79yMqgFTKxh2ct9y00BFYkPMdzAr
p1aZMiTBV3P9aMYieeKBm59iKNXSV6pOEEvdDnqCm9c1LT0b3kYfueatZE6N3OT5
IUkv+gZrlvyheT4h/U/87dXgcULNiDj3Ecpj+QK05Lwu0JBfMNmRP/BrdocGg4ux
T7oOq5uDeN8ysiQ0fuCsUaLFnJsYcevKXX1LNCrN9lVDRnha4kYJBbP2BPU/5gHx
yWYkClug9qU/crRkhdKyjCxT7BmUp7hFCKMQK3pBcuJKJ2RU7nZKGTINL7UfrHDv
ouu3XhE47wTUkTRQUqb9U3rqb+HtaJyz0Hq/fW8BK2Jt7miI747Lt5arMp7GqqbM
3MIDkshORdwlD2b0/P3U33VLEzAwPeJiu6Znyz2IPC9CJ5OlqNojOplVxPdjiq6W
gBlkiStDjvmIQLJcSKnKPjEFPG6ThSQGsMZEpX+AzW3ark+bajQFIyEBaZnkR/eb
uoH5z7QMoXUwDbew9srXWvtozPd1LHQftX4dq9zMD+PaCVRhtDnue4GDqnhsezQr
WXArhhMuUStnNjCufp/TIIakraksJnB5LpBRNGRr45ks38gqWKaUvl7RSkBLgYXy
sF3lW+av8gOZIzZPRXZfkqcjATt15uAuK23rooAUEg9qXjmloLsrhVVUC3lj4evV
/ulK51S5xxsA7SYC1MvfiZhTiQ+DdWWpGPRIy3BhAxTQnMK+/ZrrynjpIiUAJNV2
X2LmF4OvVFE4PUdzQf0IZWFINs2767N7m5C3+7D7oZvSpsB8CW0sDKwtN0rC2V7C
vkrbFbIJo2ZflBatBe3bvlEnUCvTaDPgCUJh+ObnGZgpYdWEPUO207fFMqesjytQ
49mLO1rbpZtqdzpeV2HCkFflFFoEmd7Zz9P8nrwZALka0FfAd+sH7yi8wGErbiiY
XSsqrKrjPeh/NLSRCKzqgAr7yzBCVjIk0E8OF+P47I6uym4YcN/Lvi3Id/bZnhJX
zCcpC3jC8021v5yrlwiEYhJQTVUmZ1lorG0TRXWMX4n6T54p5i337DlxJq911Hh2
WeR8KWvmQ52PIVrxC48YKTzX1+k7LmOg50ozYnwWDGNjk1cYEtLhp8UV0vnxGHl/
L6LOzPvpG65xtmM7KrbgCMarHCCtYY/FQ8BBp5zpstqQ+WOMNCM4xBDxr20iPV81
WEvR/qlfRQltMp2Z+oPTREcc+lfHp3TEfm5F2YLTILkpsvXL5mhK72Wgy3i9Gt6K
WrdgA8WPDl3epUXLOkElQYpFbZUeGPamc7TKqsWb4JNUEteCHux8va2piuvpe0cU
+kQd7L2CVUT1zAPgDWveFZGqdj6AJecTkxmWi/VWmQN9V1JmqfAzbgZyZeNNZUo7
LTTi6Yd64Ad7ebzTlDb9N4al4H/B0qRWl1yIWV6JP15Xncz3dLA7A1vmuxEZWErY
hghT0Na4unZs4wsjhUbmSCh9fp36Vg/4tVUS6QDfOdrUCSv92cGfokCFd92C+unI
0XGuLDgWGmEiyFO4WhWMMF9+agf1gStEHjJfzJIHpizO9Dp4KXYtO2jcUzhiTLvi
+lpdJY0xys278wSl/mUU2esITDz1QCPTQh36VUclK1zhPfsOVDjOAvGo4qyIaqoa
Sl8D1YtK7yrfX8OWt9Qu88uW+iIhBbXACsZ7en86GFDJpKolesC+F+5WdOmbBKAe
eDr6lPXIv+0FYZAYhPAtepMZvPlriCRkF630clg13wnRxieXeBGsr6yBTQ5POVUT
CU5wui0LVjJmMebzxgCabem4KMxN+xp/j4F+XCu3Lo3+dRugZHRy4zZTrgyWw/LF
EckFWjTqnHixvbBsL6oV2Cjdp/3ujqk+VdoAgkkxFj8HWvG7TIhhQEvtcuSqQXvc
R4xKVpHkD/5NqERD5V8I6p65kRVNgJXwID67nzGut4JCl+2jeAorwHlBmm8G3pDl
75EXTY4atzRz78WDNudBSbv4g/jAcZrP2+gcv2FZ6lOJvjVuw4MIXd/RDHDj9HYI
u24Lrw3T5Dhk6B4zeVqSbm2ptsSP0BMy9DZy/teO94vSHEHEF9MGrMv0p/GSCXZo
Dx1KcjdkI2pbeEBJ69ignCxu7it3aghO5xPfIJB2B/O+TlBNNGkwQJ5fy/6brBxa
ILC23LbfsPeWdbFhLyCoq4pydqAdoYVZA59+5EzcqLWyWXWEBv4GJMEG8BUUV6rY
hw2sY8I9uVWru31khdFB92v4yd6mlYKovQOO3202CSC+0itM1R/vXSoaO8ioyWDn
qjN+x4UjvwsIcA3wRKzSSSZI5igRECx8nQVU4oFUuwbjATbJGfuJd/AzVy66ydDo
kD8RoTvnZxI873O6ZjlzZ72jfb3mcqOdP1mdiZOMNp8tNIvtoC1ES8hqkeZ8AHVk
na3lA0vfJY89np6QWtQzeqBaDk1eSQRPoAnFrHjhBdZ4GiQl4Yj6PzVXYvl136hd
QfmhVnGx2dyqYcJUPqbSr+tWNYg+Hg7adtJnTw/apoWyq9t69EcGmVryCd1ETdKI
uqHI0in83YemBvsVyQxMVp8MHHE8xpEOq/P1zoGSr1HrGxsoSvy9NFb6XbP2n4rM
Jqdr2X1oYlHrp+4DQhF2xuJ1LojGXk33teHoKBZenM8Z6LEiQNSbTW6EPeqv2QRd
aHfO/jyjmNx+1lV/lrA3GmANoYFZ6b6HDRC4ageLCHAckj6uB11EOY2YT1rJL1YB
6secsQVCgNGqhMlTyiaiVAhhSUpX+WrFbKZ7GtKIMv76EQzQDf4MDsNYmh1UCC6G
ZkAvz7ayyrSsr6n0gLRlM5WuDwkWZByG4SuW/qIaVa9r47qjrmIOed74b2QDrzEo
RxE7k+RSJufUKCkJhmkLGrjGWhCicIts2mU1FpSmf60JQK/kL/Yn2y05fhN3oedZ
GKL7rj3eWIPlG5lqbAOgciO04meaRJ84ICuCl1WK0vcyNYggO6tao4CUku8Pp+Ry
zSqwPnLYHaUQvzkq2tthEdsPTjvyjHsWuyTpxmdnwSUpjip4SVPBotSqO7ScDueJ
AQemUMe8TWJnd9vDQvZJ2HrPxIB2umvaRC+C66ZahNXuPKJXFOPKrIsmYVBdWmTE
LDVmbtVuRnIiUI5UZaVF5ohsNJeGa5x3jDUlpADgBE1NrJK8yu8btin7CdcaOBGp
MpIIMb5/B6f25Jq+krBFtctdeqeavQemnPW6/Nee23ziL9vWjjPOhfwQLLEl6EeE
CUPUWbpWBsvaS77zMVv9WyvVByQc5hLwWhNQsvAAfGvamfKzI7PgC2gaaa0TE7a+
fxVFBGifLav5wwe9zgyvcnoCDykU8piqGO4PqjpcaHsIMbdHaGkrY+a3JfdDfXEL
sqqoy/lHEtz7wSNyXX0aBWJ24V45BLDbYhpLQx9Nv3EDC4+QUIjJ9GEFlFqBDqlC
CVzX738yKj3eQ7fjA1ikYr9U9630xEgb2qJZjuSB3x7BqXEH/2WWzadZaunGUKGT
PzfM1ZQYD8PtRBjiCio4tW+NVcIZBbZ/obB5MpKOVIyyQznLw/aA3mPj/T3+0gMb
4c+CVBYWKGRA8TkKXOFrpHLYsnAHP3RN1+EYh3Zu44Paf1n23F/aeHYU5NgYRuGc
RKcMc2CVeENKw+wgx5FZLJGP9yeQ6wijdt4EAeo9ZHNnKoBtQFa/lTgn8cAs0obh
djluOG1juf0iNN32lS6gxA0vfMP2Z2OzyxXrZmva4daLbzbBZFDUTrPmiLYnZhCI
FrBKK3nRK48VVhn68xa7gm2tHDLzzmoRbtyf3GHBq6+6xSlvNE62gMIJVPIDW4pC
6495ncEpljPWAzoqR8gpj18Z9m84UL3oUEyr/5IlWQ4SdKiLYoEel2C2Kbb8JWEF
5Nv0zDbP22y0EylREmJdFytWCk+cyzWdWys2PySbKbL/AaUBEw0L4mct6+W7m8mz
ndIWnunoHO6HiNvYmmUORGd30WobBTjOJjPIYoaz6O0Tu0LDaNwG3foapPciOFGU
0iIYHhtoGXrNUeLCZ3ajFMEPID8LKWORWcLQM9spEFJNsa4TrpKhSAfBSpD+yTKC
4uLaIgsq0gtnlmjlWQRNp7Pw0ANlSfgF4Vc0gyHy79hdnRHF2+cN6QXi6dp1QrsD
0puSVexvIvOYrCbAMX0JaXwVA9Jg3KSTRQDN9Zw7VDR+LNLAAdPDAJ4tkp0fLN0g
eAUw1dMsS/5OElRREErlTh+zOP8omhNCmRp0OhA96+D/I+kRFSU7ciZoCGarCLuX
6udw3AzV5TvoCB9pYXUJqU6TcvTIyypv8m0UE4rJykx5/2cxXU1L/RgNer3chNRc
H0NQEvdQ4I9o9In1asBFHQg7sLlC+In36a+jEUJj7ABWEEC43TGzNqb58nWvwTMO
k9JqIoEiJbpCeG42OxeNmwUBoZATwGJPC6BJ/zihjA9uKaRiJvVoSbDf7Z+YE9j1
atB/wFbWM4xDKtIHbNTeP8SY+635B2UleApNA2OUnJ+XSBwTJNIqxv3mnj+BUNRY
J8EVLFLhor7fcO4kDIFYFiDmxypCcErVHVHdBRaEUsMqW4UZSxrMjH4lW0HUVdl8
kN5TGhKZ+A4Ve/RC6JEcV8sYeAo+3cohv0ygid/P0cAhg8ap6Bu0edk6AMJgK3UC
wHFtzRiYqzmnRqnT9Hp+XrQCTGdgFIqBEcySG403tjWL+V+ge8p3nAshj8cPN3a6
PagbiX+7Tkb5VMEcZTHden8s2s3C9/pL88rfqDRzuVLQBIkAMpzEHA89N45Yl0PH
8Yh0qOrcJO/MYyLw6oufbnxcjT+JQIOzwY+W2GZfUwatF3wxJ81OQcSzISQs56qw
niuIRaCNUjdg2wOc+az/PCvvTX10vA9S39RGPXHliZ3aNN7TqAckrsIOWhWB9699
r2/H4impr12em+DrQ3NfZCFTQpx5CgOeeO6y4BeBNOLc2/zpGpUKwuljIxLbLBQP
M3YHJMaGFwxwkXwUV7uqbK89tkP3oGIkwkY2MDnJIDj9tRla3lm5aKZrtrG6YBRC
ut5tdySzfWWzPbuul9M59MldqH9S2LQiv8bmpOsyc4h0MgEEYlTaN5bTEkn6wAss
i9bkmX6bATM/hsXAz4DkpnCG1YlU/Q871fIfhlRe+9Z1LSigEDhKigLEOuxOPYv/
cZTXjm08Ty9NWGpV0W9EZRNxyqxNiCIWmzIIXSZj9++qt2Pj94uC9lmQTSbo0wOh
IHLNMNntwGWbuaY0i80kLUnQjY8V5ZrGv2+UaEkmn86oaU67ZKakkXys0OgoPsvL
EJMowz+UTDKZNtTRnbaF2AWK0lswDbWmyGVVnMQ7vBIaNTTaGEX6ULBQUE3kYv3m
5NstHR4Ij1cPZ+p+jwxhf45LjG6hEZZq1H9iqtPV++77MZJNWYbMXc5209Oxj6xF
1/38jVWWKUMbYtyCb6Lpf9dbgc4ShF125jEzNdMN2V/ygf/CmAneikn8dZAL4bk6
8OBV0m7xxNsyRaKjqhkYxaSTGiy4UkKo2giIiSCrtG797eXRlMqAzY+TehYEjUgn
3CueoZG4s1d7DZBh4PKhrWXDgPU2JcV5CvCzm3H+bHPVYPaeKqPQKcnayIzhcsA4
TLy8dxkSD6LLfwxcLTDKIvb3N4x8PsSX0NTleXNsyoKGQQbwSNxS+m9l7xKQcZVZ
hNhTSxgWjxdRWLl6Fj/lDJ1klFvJpdV+2dih1XREKJmana6HMVCGZcr/Ps5HyCqJ
k7G4jI133HDr79xjx95TbTybTRCf9MMSFlAr8pq/z2QhbDxJ4ffh7XM5UtGEArK2
Ymf4uHBUgLOc36DjnLRm/0kU3ldG8NKh8Z6BBV9MTK7OS7T8xiHQuggTjyXwpAkS
db9UsM9NbErv96DmF1dF5g9hc87nNB6ykf3BxEigOZ3ErtmLf5AAW+T3s/segBIh
+w5VczDhaGUAEv1p5LAzv6Zm2l+6oMB4BgHkao4dBiKtCTQ9OTdPsV1HlTN5wWGi
5zLLpScfyyyLSpveeiM4rgykiZ4lz4zdXuYPg3fU9oKROGpIsSJlJuoiD3wvP5uG
kUM5X3hlFzskkA/0P4P4i3B9KNVBOdYyHY/OX+Jw+Q6aul9mMECdfR2VdM8p4jVe
U3UVRVYHa8FMBcaWTNLGRSKoSgHFqNuoxkYZpVcz+h8stUKz/nboiZMs4Y1gxrXk
t4CHXDwAmmdV+bZuyoPATvjUWqPaTrklBAVjjUzX+iJ4QnVNihNyXYRia09bH/t5
KTqxgd1Cf/oU88EWIw5K0W/7gCbZDOBMwzuWGdY4FGOZtA1uFzIT1IDMaPluM9ga
RGNMx+KunEvfAtSnaWvhgbX85FvZ8zuSBSQC+uKIgXOdhok+wULGKbHldSGKynBA
uV1i83PpfyPP00IBXtW3q4NNYX/dTwrvq+ByY1W/iTgRx+9/H1rRUIUzNLJWXSqU
ax44s8O/TqhlGwOb3Q0iABY5bSKsJ1LsmngsLhsabl0fxF2crjcmzJTTkNhnX92H
PrTtlMKq2yLZLeYzFRXkmSlosjEEVoJ09k9ozs6dDK8TKbLZVgQWtpiUzfOIp26D
elyxNdOSX7smMlsdP7Pt0npvqKyBBiW9LWfgFjTb5MRrv+ljyXu+wP/ZEx4BJiL1
V+qiIHvSuw9BVsUeKmA++O7kB1K1wLuZyNsVsqZu9RKZaRia5aq7k3lNbxSGtA8z
WQeINBwzPPJ1Opl1Pu9veIC4irCzmc0wZp86k9FOvKU0snzMn2+C85LmCadKDcRJ
F8LFe+6TMAesxMfY79ioyCNUxVcOuM/zXfFHEZFyxKQx2BRUdmsSThHC0kZWIS6e
3VdKjnjc95VMaZygDUiIbFIbJ3j+4SBU99ALvuR9oXiLIYlMgAsCgWbMWZ9Z0vO1
Vpm/I0ZQN8sApsZyuhhLBmUxbX2m3XlztCglAmdEjzp7u9qa3kLr8CFQ/4MYHGmn
0Cpap3V9PCoAug7gZPfrPz42BTl0zNDJPgJghv66HgfKhJjS8ohPjno1NUFJcYf/
YTe8KdHyWTySOqjS/eeeW2VQDI6/q1QtBYukBasYxQYbjiz90FVRTZ9Mx8ITKZjt
NDTxfYmLuKEPT8gouCC0eLpYlxJbdT2CKboDxKKT6HXdCOJ0A6pbNuUzGqGE5NUx
G3pl+lKLXuqhDiSFM+L21V9jiRiBk7tT3QDL0AbOcF8FcFCPzUhGoE585PqQh1q6
vgcTeH1do+ulkangeHBdLHqK/oqzyQRxaZzdizprI77lsPWVj9IrJnxUTkhM+asN
1iuTYgglKdOqm7nEWoKUG6LNsC0ZoFSNlws/4GmFcuvxD7pm12YRsKSAkHyJq7Y0
iLyfhSDhHN0s3FUMd/+lH7mbGAJQ6ftNEWt30II9WGArq4ZYjq9VOLhoeOIyzxvU
y/1PAD/PIY0CGon6syycNXk0FSjMUB9yykDifYhl78pGNgny/5AIbs2/2X40BCiR
dfOqy10hoT1DxfjchCuwMNfOeUh5q4wmLf4jOqqjTgpltbZKNXRTqQP5HgaNut3l
pjJt6g2AjNocloFBzEfDjgsPoA5HsW/wVnH6x66canjO5vUX2YBuCL5iTyNwJaiB
FrXMgS6+dCSLZ92T0+4LKiNMCV3hCe9kaLqUxHLDlhj6hHVQ9ETt3cuZ4SqHs0kq
2itvxCrHnfU2i1A+iuAXbN/omOgrmwQplfWaGhuAM8C/moPayVweIicg0/BBfJ2f
kJ9po5sLaCjTwv86WJw5OI9ds2t/jNCu8r+pn441lEKjAPAiq0bHSc1pYE2Nal1p
q1vV+PcD33Cv5f8Qt5Dt5nKuKeMonl7Z5f0/v6lJpGgyJxWgnKhXSHmQyKe2VM6r
/VyNUZ3NkTG+ROBaJBBCV7n9Khjs1mBx7OWWihGuhrQA8HyGXugCBHV/0kmrl9IA
td83byAq2gA71VcGGYRXsQ6VT+6i9R5lLYceJp+/ZV8mT5EF19uGkWtGkdHxPVnc
Qrh+VUM6RdNdbL5uBrXXJc8z1aTnRFlvzWMg1/dYu/833WDLpPIbMROGZwceg44x
1BW/7YUNXskUf4ATCCzMuDqkI8c2/vctiNlFPKxldoV27PgtneZkIo1eqcnV0AkY
IJpGpGki8NDdxbQtqZQEtqueN82U3rMT48B5ufK6NzVOgh9YIwa8ZCwK2rHk7M3z
WdqqYkidVs1Ve7SkN93+QF/nVJX/M/R0xgvRDWxZjYyGFRsDuctNT0XV974S7U0N
B26srdmL4hu89CspF8reYI5TByPliQCrgkWLPgR3r9UxpdM6eZ8r8fcnUUaR1Its
G9omCqmphhh/H4Fs16jA6wTmzrzl0YvQCAzQHzqndIlYLDTkszA2YgHSVXjsHpHz
9Y5HVCN6+NoaJslvJLi1H11w02phywaHgJv3+SDehrKo8oRt0nPcNKmyy2U0cQE2
mT8gG+MR5TPijf0ZnbMs87p4AsMC/s+zoSjSfUeFF97YOshCLD2diC2roZuC5MaC
fUqE8KemZvrN/R3vUI7bEScQ29umh2F6f4x6Ah7AQ5bm0Or+zSXtYU59+2LjOeA5
rNRf/Oo6rTvuOan6sKaboE8nMnDiCNOhac1xH7ByZkBKKgg3zOUarmu/ccRTxh92
uNyzkNL/+pntQ6Er5Ti2VkeYOHGK0eg6AzWrMF/JArAK9X490UVgBAyI6+j1EjA5
9LK1eJ2CMeNIen/bgxhg3/cQgJxh9zmjSt0FKIq7SbFqUAg9cs5pPm+ch/0bbE0D
g0yt4U1fVB8yXkql+yJ/oHLI1Zzx5ZmEm3oJmY6Dxjgd3zSVgJbJnf8cn+9+kZTX
41v1ZtwRBBaQG46NDI0mxmAQtHTpk+uUAPa/Rzibwme/NywG8XVpGAAtL0NoibEt
PXjCKg6wKKlGeelGyDacFHBw2FBFpBPtUKnI59Z1ZuQbwvjAElW3pAmQ2rszLucv
nvj1q+OV4WsxyP708Vrgd9uJYLmCqRgnq0KLcd1QziXtFCTcICzaVEbP1pwfRG55
IDT02HA8U82Ek08TFowUQBXa7byO0Q0rBkTVmvZEKn8eF3FBarOKlJhcmjlb7wZu
aie/KZpu7QgawckNKNaDWbKIOE7bNrvswFDCmv7eXpoKSkKQlFDMdzCj1AuvLa/c
QqrvqzMHEEbiv3YbjLCbujtDo3pcr6thUU9x1yg4EXKSxSLRxwSMX6Ou+lYSy+8Z
M1eFTkr0hJNqspIztsojeU0JFKjqJv87DXln15oansf/eQambJZXzpaV6BZR+zkk
KeXNRxWVfro3/WbU3Wt+k3iFOAkRKQHFLCVVHKyhq6qji29AqdJY9Fj0ajzTgeqw
kv1GAR2GfJQME6purg6RN6zwGw8BmCt8GI2qEXwkxVvBo0iO4DRu2H0Y9B27wM2Q
jGisWgs14lQXgQErewMOZEQzvnq2k+pgNkeuXZ+zkqlOiO+kHpp7cCU7WjG6/QlG
SM0T913jC8O7moShhkjE5oYF/xniDu8Bw/WL8vnLgHTpPeWDKdYP6xLpXbwKF0GA
Q39W6IJlG0q+3sxwG6BlZ/MVtPwuTfgJbg3+s2iKPhqF77uuC/Dc6DBAFwZebnYF
rZ+rNXNzs2iQ//NpgMVPh5gAuDIqu03fGa93PABjQda08iEyLX9xtMk7jJLHx79Y
oOWGQOprV6KlTWTJQFBbQf9UDOomUKRDAsNgBAmhJ4LHAiQQe8aUmPndwINNT/Nr
OZ88GkmO74dwDGDbmcAaWUcjrxrlsLbbcsHTLdYNxA3lZ7QOGeTSIPLiLufsipki
KRTh+pJtYEL+4omlDsjglN25KUgEoyAmBRur3dO8/J+qYc93hPwsCpqUx+51dtIh
RAa3vuBTjbDoFPKLi+xNHohxutHVfTaVgDYigdomDZnQmGZRggmTpEm1uqyt0dXs
sWOCP9OYd0njWkYVoYEgScZecVJScx0LV//qsE9OcEzPnH31O/o9LVjCJoQaTo+Y
kJrJrgmFdeUsH2JDf2KdaJMm0LbFxWdaZl3LBp0hicwKZXm7HwxDesgMbNz7i3OV
692rrAN062/aWFlkB/PX/GB+JUnKUk8tvzmzUFtV8FeJ0oWSuRdeNZVtdjgJKAzk
nR2TnVc5XPpRakXiWAZH/WH4kkT4lX2t38V11Zaol66WEpPBTybue+WnNGXv1eY4
pkteoyPUgymMIWXnMsj1uBrz27xqkyHUWWUAV332/6iAyIlFsDi3/c7I2/Qz7WNs
oe25Fdm1wosjeJfyzWcKoVQKW9TptwZeV+Rn706iazW+Q6cao9dwrnr8vzHSrtUs
1cU7OxJWWiLHvICduV9HFOSaYA6mHMvs1G5Jn52+iKPj1lXJ+RlB2rs8CRrPubqh
aD30NpD4Dbjz1ZNpr8QXtz8FlPmnLAOTANC4WThh2Xd6cOhAjPk6URmS90XCvhNF
MH200ma4YqqJl4fdrRnq4HVqycpgphQWRkrKNIdCIhf1aSDeTBa0V19JRfCGBEOM
+CIjGdiiVCuHlpQr8jnyKjWwJxyRB+RJIswuqUNQubgU1/j776Jht5lxi6KtB9V+
aOO1v+xaJmiSecJxzKbX5m6NXmIwv/v1wjHnzk3jr1MXsg5ySuaTWoRL2iMHw4ZL
WRHxBf2Ga5g5T9IfcuUj37NKIDBjZfFVE0kLoK21gSWR7rQ9xI1K66HXn7Je5e29
+lagYvbSi4OcqqsGZ50kvf137OUuNhtJsmzS6ypik7nqFslmnlexiniveSRIS2Hc
6FziIi9pyKhmqp7PZjbZFqwj/68R/ZSy2izOsjKl+JWek9uvi9UQzVWQ7f79e80v
ysdhS1DSpPQlp/6nyg/RaY/jjtpwaTj20MBmIr47khmct1GuIDCEehScC3Z4Hf46
6VCJK+1ARnMzxxoNMyctyPzw6JddsMomazrpEHlMIZHN9jypibpIQPtc7HPEbJw4
fjxtsoPM5O5Z4oHmsqFrv7oPAI2+BhIpv5Qf6RguzTprDvQdpm6V30W5UZ4AFdGQ
kaSC6mLS0otGKVUOpHxTLEAqGV78stPJ9sjWo3gVbKcUFbjTqRClQBkpVlkXqtdq
UHDKdc2Vqm5KVRx0UGH4Yp34NS0okG7lYNOXSTnYcjSntR0ZWNn0HhgI/ula3RyD
T8afddg1HDLphwhyzWzjgu4vhxf/JUV81+AIHg9PFmyLGsRPrj4MC1e4pOEXHOeS
NrTviRYyhtp35x4N5oRqQkbw1qsSfPO7Ht3lUu3elNC9xd1tHTKuWHUtIw4VoSv3
Jm67g24hVQb6ToUU5cuGZZHcxEdPuIG22yybcPLKXAuV7XTC5IxHsCDJgIl7ZkG6
5tCfO0yUBFrHzKVPcXIVbjVOIcBfRhW0096NL8ZMvvWW5UBntjqx39EQXeI2fU/3
Rf/8rowPqQJ5jQfMM1IfxqjX7LrUA+GIl5sprX8M712xb+kj8vq3LjyiqnyW9ykk
ROS0iuK2nz1Qn83+E4oeimFjbijtnVe/fw6jXN9OJfhIRflIkxU7TTMql5KUtoGM
Vc48c1YVFzCzu1Aq1foshoEceXux8WPjJVNORgfA0V7HTUbAD+T0Iktzb6L82wHo
6MDf6cIxfIPv0eEyva8muX+lvWOZhPTbCt9l0k72xE1taMW0RFNyOTtOI0R1jg+d
D9j8A0HuQyvN8CJaN/qiBdlMeT7oma4DikYes8sjhEFZKuqfWbrDCQaJ8Uj9Ei/X
Rpqh3soTiGhXXd1hbBmIdsQ+rN9cOoglmILLodvbhjI1/C9HPS6W66xJ6nGz0AlA
83JxNDImG6ZXgqP6Fa4fiPBI68w19S3NATFr1u08q7AX742BoYT7WMLPaseG44lS
MwfwHi17+VlVWUKXpRQR3CYnnaTwLht1wz52L3cWbTBj95/LaX5u6GGyiXX630ab
Sw4OER8wnr0KO/uYKPuUCx85ASCUNaT9ArALF+S+c9G0bm5hymJJnVXgDwIEg6+O
4NkX+gYRlO8n8y3I0JtOofFq/w45TrEZEgOflWElEUHwZG8UDdcsxx9xo3jp8ktX
XQwJw7SxZkziH/WzQpxmnaZo4D8FtSw/H/3wLeZgjJPlUGdPaIRE2J1wp0exdXpU
JHEqBY2kspxEYENC1P4PgJ2oboK2IWNSX5tKfF4Bf872aM39bkpMNiGi6UDPe5wt
8X/xvX6QVJLMazas/aXQtQg2JP5Ec5RAz+kDqlkfwdlJ9ETJRMTBrggBp+wo+eC2
kwcOrbKor43s0ku6PKwBCAR09BU7sMfmzlNCZO4fZrnbMX8Ruf/0EGzr1DxtwIGX
y5BaLIZkUphy7kLooOeoQmp651bWen5YHIlcPEEKG5bATsrRI156aGCrSCsJGOLE
OHjHJX/hq+vOnpIrw5tUijVppnX+pPGXcs8yIhJAsGbhIExO5tJDR/SlugBMDUDn
uCuca3nO0jQyq+74G09fZRHwPspjP+ud56OABXR7q4koMZuK+ZNuKPOAHw2j6/+T
HUK2wgwZFZM4Y90q83jGPiJN7uGmt83/nlys0AbgTuYP8kg26VQswfPe6CksCy7L
bAB6KUgaYMDjK0jv8RgAHHjZ1/5wqzrFzXbO9UYBbv1U3YRXkoG9ug4kSuNFvb6t
E0CAHs91otveMeGvBZLLTovGDJDrSRhpIsMmlmgaIwAVX97A2QFgjVfksMbNNzWh
ajMwaoArj6YwUGQRPzy6jkrU4SEzvb2BwV9tIx/pdxfIaxs6+kCPI+vJrgace1za
WIJHmC5DIbVe0hLgKSTGUyDK9wcuxBHEMqtUNMzd4iKaw+7vcmpu5Q/99ts9I89s
Ih0bjSUmxARg2W2OtQXP6xV9WXCLzMuIo3nXopJnAUlD4/PIRR3Wd+T2h+67ZfKz
0h8DVd7vE/MqLM2Ia1zyTZFJlE3dUnKGvfZF7zVgt/8JDnAR2aZATYxQQqJTTYCn
mpXiznFU4FNuAUtLhXtdwAfk5D8afkHY4sUQJKfVC6HKT4xRb8E9AeCpWbEYzuLO
BppqilvXBlzCbQe4/i+BmrQAJfQ88PnbP9ddcWWFGJ8JK4jsfxMe99lrOWoXgfoF
kNSFxLMJVnVziwJgl4tTB926+YkoOFOGQc2Xx6qHIxo6MG5Noabkok9CS2Ug4k7l
d/5l8yNCPDwHSjkKBLc9zVFsndw2RN5QvzK6XJirSk1VGa3jkHavhxbkRDPri/jK
+9vC31slIMDRbZsrFylvocsTNyQOvAWxqLU5T7EzZqPKvw16pp4qhCCeZQJ0oGzQ
/DH2Q1SVRAqz8W32r7dr9UXOemZfLv1pRK1E5K59UIjQhmZ1tAsQtDjKt1rceuEX
NwzpGH3qI+p9Wa8lDDSxi9OOQ4T9aGnyA9VYiwbm16LXq9hmxmQnngRKjcfLMPHl
uKqXk3AmK/L0C0Dm1eVFPBLqV2NevRGGbKQDzlgG7utnlVLZ+Rf6hPOs9enYMWsI
l2iCNDGOdB6rcDr8k9MXH6H8rvTsD8nF2fa6r4TD9cTd+ORkHds7wZ7/u4zjz8uG
oN6/PZDoKWEmCGZ7Smy4YaI44U2jk4xQFy+hEOI/AmsUynDbxlpMDpzeMaStgKZ5
xz/wXUv3c2eaeqnSJnas/iZ6LGG54LmqFdz8CmJkeFdpDtNqAlBK6sYF1C5N8I9+
RS53f1HKhV3wezDX9lPvfrmIiN88ZpRQ/w+invDtMBHzOoxeFDtKxbm/8A8T9Vfx
XywNj3AE4Uqf7fKyVGnJzUDWsbPc0/RE6vBmE0VoHFzhnl5k0rfTs4M5FQ+K5DEm
ozsOgSG7glG8QIJHK4AOtNurlygwVJ2/ubjL6Lq4i/7r7gYPnVsGqUwFxeFW4wn8
tZsaeyCxYs/O2KUnlCUpn+suDVUKE79u8cvVtC5kMAauRYJ/z84huPGpJwCp8SPo
nyaza3veWdTHaZ54SFcX2vr8+v7daepiqUn9DddPysAfCP5TcHl0cxLnq/O5gzK/
Uz7NL2lRhaTWQbR+uBizPxdOcC+Dc0YMmVVMaDS/3nJvKIIcx1nmffcENQR+I+2D
uddy0CRRyB4ltrskl9h9WOE8I75TFHHHQeJZ9LU9EQOK/UGVl9ShJaXL9s8rQGJX
u2euz43cJoIVWj9LMbQpqCwrMye8tqsvcbTG5t/D64TYJKtSFELGB75/rDv2L3H8
lGmPnwCzg2PHm+/2gv9PTY9isQstLMFvdnZZTTZCHv+/wAb3MXy+Q0yKqFNTqPGL
9ooewM3/2OKfCAGO31sN2klanrb44/obPXC46JUi6hfDh1g4N6k9vcCjBf2xnd9x
4XJNjxe3KDAFpIk+0Wm3TYcDDoHIITT/+x/g+/n9swpKg1yxcDc3/jnDLCfVKcxH
CFQIRuC+urvLdtIhc/EM5L9ZOuQsDvwqs7UFSz8NgLUebNdTHW4iR7NLwGr1JEFt
vtbWZKR+OCTj9XZ/dImJ0oWvx50mF7eWT2sb/ako53pcOg129+3FMaMBTsj1fXVl
CvFu33y2XlV0GZmGy+Ebdu8c+Qw0hRc3uVqrOquZTu1m4hNSJ3nt+byh3NQMoaJB
iR+V+TPO9zZPK5HreEG2OMoZTAzx0ah5e9vklGSvyFfGKxv4wY7A3bE7kGO0ADA9
kl0GZJb2MtF0e/OU6mE9/kMRFnD6Z4Q8lZKFKGNphD8AX2lcGkQPAaVa3Sq6bLX6
+m4iXYlr2izUfdCKcK7sgnkc1F5pcLvbKYzkPRr6WY4VUX653A2MQ/YmuaBg68B1
v8VFeqNEs4TdgcgFIQntrkFrooZVfJnAmbLHDRODisA5oy1+SGDJk4KVwycgenh7
KVtx/moOG26HsBArrerN9pThmNmWwaCO8At5faNSesUhO6/7oKTJP1Hja4t1ANjJ
SazAEgx5M7wScmT8pa6A7OaPsWME6Tkvj50pelJuuXLJ0tesn4l7D0buQwxCbBao
jpFJ64lgzokmIHKVTpNOF8Tbt0mg0d62mgGXamuMHahTgXogr75ZG8RCxUL4+gHp
d1x7QHkzRpLafV7UKMFpB/fjsUVGvKn1KUHrI70syN0NQX2yMP9Wi13uWmqMnklU
1MpOUhHEd4KAdx/+QPgtR3eMHixy0uybf5zSKwAYI3SInMyAVTSjMbRzbvmQyWsP
cIRtVEWCdb6GXOYr3NVYfQJxELtSOkmGR2SWm2rmAbejfblHsWtzOnkjkyVGeV1c
U2ko56+54hw8YYODEXwVxr8DBl2USYj250mOtTJRz48Zy6L6xHCYbLVfs7TXKHGE
ofivgNrbAe1x4Orq5NknnrU5I8fNT05rIQakzYO6BMXmMONxHFSrOlUz+Y516w35
38COIwFzMSBR8BQWNgcMdBJiS+F6AhP+Hq/CVazpgCAfC+N7x/5YoDUeD29peKN1
5gdQu1x2thX1AgHCNsv+x9jcuXG0/RM6yDuFnm0xjxQ5dhqSiNPMLKd82Y0q3X5N
vt6aloFw0zt9m+G6APaum+KZXIVX1A8PPh6+KIOabU0n433/wdZHB7OWiDW6riFJ
yazw2ibu0Smd7KkWl448nE17McIi4TJ4fkyumh9Cw4pHl8FBPvy7WrQI7TB7jKhK
`pragma protect end_protected
