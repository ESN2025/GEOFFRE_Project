// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:25:51 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l3YP/ntm2VEVvmgKR3q1aTb7/OV8phVfpHxyA8uhs/YwDLBJbxQ3FyQY5nqGRIWm
uoPNe08O7c8/9YkP4/z3EQ7LNUczU4Dvtrao5gG678ZuiojRkdTYXbGGZ+e+ZUqo
j3G9CBTnz4llRNlof0FbVtsW0fjRoaMdIPvnaZ7DhLU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14992)
bPJXOcxnjQ4t7EpyH1pEQs41FyZf0cTRDFTDIK5fX/Db8OYyif0L35G2Z6qaNLt4
A3Nxrw9ySdrxKdsfOs6PxbkhhfnLEwsdjLwiFDQPXe6ApO6UQThPHvi63ruE26WR
tccqqYC+zPnQMH+ZohRrUT/IPga6nsrkSw0PMyFX6Yp0Bpz4x3ROVg3VeGd1L+uB
PlleyxZD13nOfJB9xL/DyqGsHr8xdOOpc7qBMSt7IcUnf1vBnlkfaP64GmZ6mPSo
z1mTneTbJ/lJm2RidJjuiJQq/utBfB6GPLYU1FPN2C0CZ5ZedPIAUP8sJ0znSMNg
H45Q/W6YBG9ViZ1t2FMSkxCHycJSuQPYrBdkro4YfrJ66GcEwP8SrhMoNyx/tZw0
x9/IIgZOsOzPXx73JsJjAlXycj7BDrHmICyk+dQZFisQJQe4opnkLYeCylA4iEFe
JMTEawXZWt41yCqj2C7wbzAaQOLjuFVErH1AzANi8Mc7/MfNMI68A0xGaAtQFotZ
vKx3jCNj+znV2SOASaQZZxFBClYxpthe2aE2qnhIuqUiLp4RWT9Zap9HMtwxdCPC
+hdPTKcZAcUKBxzNe3FfYiQgb0W7VNwqo7tgNKi9YktlL9DQI15wV6ezO/x5ufTt
gqvDT6g7k+vM4ZB3UEpN6H94ri/9hOc0u8YfrkwIJr4IaeHoy+JnhQHF93Inr3V1
K3AK8ldcRTfgxbBlL6OFP8MTRChH7Da7DG15QprI0yswzZVb6k3mXna+hl1RJ85g
9PwVrINjkomdfbdpyIgZHv65dgCo5G6TMmotulBD1WPXJJTfLQvNyvOenr+zNKUE
Bt8U5ibRK/9riuOTmo/a7hWslSzjd6g5KgTBknLCSy0S4iBf8Q2kc9kfx9LAkooi
iMSai3kL21S2XKLlUiJc/vOSIBQ1op/9zcYHhwilMHUDie17hQyL57d2tiHug6YP
vIUnO+G1TCVh9vWuERdjkPcJ7oC5MJU2ePugp/6n94Q560PRs9a3KsN59d00M8KN
8v6J0x5El5wxZj7+1ucu3ulXLFf8NrOzaljxx8t78nSI2WmsO4wNN9K56p3qDBsa
UpVSA1mKSPkcRC0JuFzYo2kB0vOI17N/R2eHAS1voj8fKFA2Gx1W4FBpRU9fLXiy
HupMRH0Pgf1GMpPqwO6u4WvTXNyjAUma932GGpSOb22b3lLyc7gItJX+nMDNmLvm
MlCxvkoOBBx7aVvGoHFY48EQV6RJHIiDboqou69QFkwX8f/V6b9t/67z3cQRzYgf
1wx39/1/REtCBeGiG7sTKjFDH69GKS5cEVqQSgtajySNdpRcQTBGiMxu3CMzpPkJ
VGhtm7jTxKmTDVihHBExmn2bNn1ZecArdSWiTV+uNHspEU5mRqNH+2eqCavQVruf
IsGbFqs0enB9vUI9GMGPdnsXgST5N6+hcPPDxBGy2V0QfewGbu5V8AUKsPzx8LIp
0eV8+HuMBzLIjYq7TuSLYwDiHDYLfSrCr18Ye1MbaXReuxzceWE85bhcVhUx/CZS
6v5nX1lKZyzN30ngnWNa+UWXMZBxp/44WRFHpSMOrOrKVPgAf1i1RbzYQ7uMm4uc
vpKtWZTJMGnqbU553fhiVKFJQGxaxmNjcFS5YbVS8+RywEs2OzeCO2Y5nmH4547t
7+jRWSz7dkDXcQcisenqOQfnKBdccMZmtz+E8u43nnCehWHGMPbnFB2s1HQc91p9
1A+rki0lrxHUP6AFXUSk+wkKAx8Iydeo2QPjPhRxxJyx61ktBM/4MNNuJazQ3s63
viHiYyqwZijZsGJza2A/n9DQTY3CQx/Ghg7V0c30UlTeXayWlHNBu5uYJx8ouX2/
9lsit3MKbpblDWNnPbtF9RETjvjBb5GA8vdZmBZS36UL7bcq0ym+D9QCqwOI71Q1
rJcny0upbcZJR0a7D3YS6yq+c2nYZEF2S+2RaxcoTPp2l2Vwsre429CaEGY2oU3C
5G9ww/8aZeCCA7tQ/3XT79iPv9UOyGPvLmNaiLcHDT55gVgDoIi013dQGDffRYth
phsHXb4R6rgLA0SYq9vPGSenrpixBjzKSAiZ/0BnxgOew0Mot9IW2MxNm7CeG8mU
lpMACby31+6mrFPhWZj53pDA5gmKXH25UjQKDH3vIwjW502Vp0p9ct1/Yew/b7AB
OdZUwrn7S79JEaockS2smABMitvpLHNF5v94xCd6wQ0qm0PmBB0mp7RhP8HPlDeA
Tv8UpXuDE2JrqF/XgnLWBTkBinttIFyqAr3q8Qq4EZ5pQzTuE0f3D1f8SD4h9jOH
UU6eaYGNd9NvsaICbDPPtlTIgLxUwXUyZnkNp5qtG11UWXJauA/wVn3N1h+fPkVq
IsCfb+ixL51FBjq8zcSwAnXNE58vyoKr3uiUaloBLXTS6lCpyHNAqbbLXE731dsf
Qs5dOSJ7BIyG0/DJ56+atw6CqOmv4azKVL8jh3SG1/gh3Smyo7+g/UiAZNRIpF+Z
pg6HouuqOSVr83v2/ZZ36FsPLLmBa01L1RJ7xnLODZzrFtgvOSI+s9qkaPQ2dZlE
h8XkJdsnaoaw1pqzHVgMX//LKUp9rKCSSZe0+DIaDQxchmHfxoyz0odEAm/hCPCx
EFogBo9EvlRSBPnV6RQVzRygXAvxPizl2ZrLCJSx2sHd7q7idPfdJFaiPa//umeW
JJUxy0d24CzHfXylx4KY7zTlWuSA+EEteB8oVWz1Mx0tJDQSqq+pyKFEXrJdzYag
Xq8JnpH6jw3HwUhk2TsXUO+WIj7IM5WUFSDBVMfuFidLNnUZzKXD5TMMfaoO9gAt
Svnaa5VcXwiKH3qHi8SoSLfMxfg4XNQxWK/b1Ds3r+ZMEO1oEoKxIvBMmrktdsP/
c2Fkn/wpA0TM54OoubF62Zubb1vTK+qcoEXWjdXhmTdTgpBYUHah7eORt1AMfKfE
MV8QQxVCJKQ9DWO3aXnFdy5uTu325eFqpr8ZuHcMoAesFv2a/ABwnYZSFswPgQzc
/pTH5jl6WOJXjF8puS3R/99xUpzutaLmxUjjXKkyiPAxBwlWNrtOf3IJfuzk1oJI
n/DhIS9Z3YeuJ2FoGCN9O4qUCwXlIgGMoaAWPgtAPxjrBhDMwCsECXrpb3+T4TYl
9q0WeL+VQyW3qkY3Xmw/txdTVH47lUlzDNBmJ/740jHipvEUmtDpUSEOXBcfJ7N+
pbx6UmqKIwpcnhKAuWInUFNa3Ah48xytmv5bcE7kWcO/GBOKfuFJghxBGlAAJNRX
GNuuYplr7MDDLumutUVbLw480oBTTsLaYIO4pSTuZRW+h86PwIz2FkpiDdcK7Lg3
9C1RMjXijRmm+0wkfr9G9utxX7+nn2RDegY0TLQx1rC01MMRwmY+Dx1YgNnmnNFS
0xl/7GFp/C3P4DxTHFs4otVYiR/G/qrsgu/RV1zm9ul/ejva/gAAQkyrdq7NzD7g
+6U+MdcfM6uEjxi2lP9e+Q8aDF0GTNxcnR2lL7yIgihQFaGtZdWda1M0S0pzdnM0
xDwwlPClnEQhyPF9/B89upu3u20VgEU2ettfY6DQ7kyGFcx+Wt7RxahYNjhRfXMx
9uA8PXCbyvWe4wRAYd5Bv8fBKgBg688us5CYybIJVfFevobPHt4r24wz1Ult6cbj
52V0B07AmiZTZ+/pPgRE2NCKSwZGhTAyuoSrATl2YUMhBv6kfFmO9Mf7aWu1Y0+g
QwiuoADaG07Mw26HueYy0kcwz/NMDQdZCavG1prwx5NuVKB0/Ssbaf6J25/sqPdl
RA79QXNU+enXDNlOUTY0+7sL9m6f0eh44vdfbh34zA+8KwuCTXOB388j46yJsOyJ
5IY3dFJetpzp7Lh3OmzAiqnw5P6wbiNzi3hgMdPzXvgv4KW+b8pBX2iZUMbZ9DL3
oCpN2IVPBUC1TSMMf3nMBS/r98ZhQnqJLuFAD3unXz/Gb+yhwx/yIqAy6u2vWwhB
geKHLf6Qms6dyv77SIfHv4u2aztpN/8d0OxfOaHxkuHRB1LmQADv4wl0drJ8zvqb
e/NYLD/ILYEJfajbuvXxWAU2F3bJPiF0nG9cTeiClhTBnFje0z2LXTBpJXOUI3l/
eqSh9HctuEeM/0P80ZxRPuZ+ZCi+94NbGRahxcYbfk5ritqwZVs91TZzOf2I6MTN
TAMdlyc0xD/pjTC7YjS0H4w2047Vt/BJaVlEcN4Q28Y2vss9o2Sgv7RTHy7sTOS+
Q84dhCK4KFLH1wwoQNVgUePurakfUWNQW4pssPqxjZqOZotPsBKB2NIey7h/NvPV
4qo+mpmowLUyGXZ4cG4YLPRWx0y3rXbnEtDht5GeuCQm4jyeVXdWhc8LYd4b9vw0
H0cvn3Rq2m7tzNIoWhDbQLFfSEApO9d0xiGs8e7WoxcLkS9rZImSsFWTRcLVmKBP
yxpxLjDstpLcAHqBXTrBfbFeCg8+my6SsvG7ZmS3kQ7aSR6isHPBewAoXs+HUJxc
DqScvwFYNndrFUeha7ffTeLpwf+JT3E6P3W5qYdFnCiU+h/Oe0G8cJHk/kpKFXzx
hpkZLH+HxyaXjo2qhwoqsSxK9H3C3zNA//pCicelq0zmZgN8Sr8LnQAgYG+h8rgY
lZwm+0kBXAiFLRg84M4412pJxSdrGmW+6yGYMwdkbzYYYzrU5R6NUdoXnTv1biNo
C0r/zSe5O/ZSy5iY7oF+H4v6G0tLZDTzaar1hEu75wXuT2JKalO1poYXtxlcWgY2
fghIxhtg4KvzoU3+UeyLKZIACc+1IOPhiQaJCGaQ8D9+Sne5kfC6FytTzCOdOkPy
WErYXDeKvt/C7VfdG8l+F2QPxUa15DDflGvuIP3uIVUiItpJQzza3JZOJCzYergY
F7ZbYbzmNzGKmE1JFs3BbpyhFVaAXiSS6omieEjoUXJuUvnd7fkuzT7mlNAd2F6d
NOHMaIv2IFeePEJyOwX6N6prh9WJQqUVuHeLcMUr5OdQoWI8quSosnLMtam6nlAO
n/gDMoZxAkcWedC3N8mHAUT/twr/hEXklf1B2b1L8uCa3aDbCOOrQA+gXowDz9R4
r70YcymlXZhvq5L8CHdkNa99qsR1419gawOfeFlQZOGYwtT6OC8z92IgRyPUibS+
p368Nhg4YWiBOgtWluo9nN9zLadftN+1BCpYgyBNncVjdV2jDU7FUL3Sq7zU8NSw
eYX1L043XNEd31SV0aWcb9RGh+ShqqFgTeNrdYEWiOrmFAtBBRtR/CYjbRuGSpUo
s4oJnZU87WZWNjFcmvArI3nh7zGLbvbZkbWkiSYUlBPH2xNsVRthSmArftDrcW2T
N2/VOaIM9sqfStHaoPGaXkFWwgWaI1ELCeVVQtHDxAONxEtHiiMO2pY7NjMJy52L
d5fbxIeLyiEcTZqmcS8DcRhwaTWb2vyrIYIg2vOzYOxJuWiPL4WxfxENYSioJki6
+tWm7gTZpbQAp9Fa7Levc3q56Ri9RLRmYQsafiBtDTFnjIqHbLV5jJwyeDC/yxfh
V2CwH+gZaf+8/nYyVkubXAv3NuiU9F/nRS+U64gWbMAE61kASdk8giX93yM4I6ai
nNm4Q2qovcAVJYCSrXxi5d6eNBiMK+TAgF43/SaBkHEV/cMmkQxIpnbH2d6cbwYn
D25PsJleIZ5csBcE8lmCr4G7g8CGB4YXh3HxfGHRmic1ux1XJuo9N5WfSCrB3h1r
T5kWigom/w0nSe6vN2n9FXTfUInM4xQ/UdDSyNzAIvH5buZf5BfV3gTVszIkYtpc
wQHQ3URQxIb4YdWK6x+YpokDle9iV/woh/cCt+Wcm0bF0xW4WQkCTwULIcTB2CfK
9Wkt0/c7QMcesnO5qSoFmRySmC5HP22R89cqzXxAoG/H/iRMwhtzFGrwfn6+Lz4T
qr5Qq697Dp82xvTyipcSyjdFPrDR279xfo8yLKjxoqa+GlK1JFbUAodbAmmF5lF5
n/XAVrxYt5axd5DWayu4NpHmJGuqqK/lJR8h4K8yTfM5lmuKfgOLsSOEgniIBDOu
kl+00pRdV2Kix+4XE+nrNEEpy4adF8rueofx5nADBOjWgdgKbyCdoqCWVfyi8IRU
5ZOikq7J0lnWIBq7FiHOE7z6votdP19LwzG5r3qqFf2zYsJmsclj1H22K6uxNKMb
CSAo2TqFitFrr8ZUc6QlQKXcrgD6M+G1gpZixwHyyhbE2VLNIG/tFg/iXHZ/Vb0J
/iY3hrbnd7gQwUgavyqm9bO8/K6kEVM7ae31gYSc4UtJu9HKoDe2S4ovvHi721Nm
VeOkTsBuKxnwpGj+gZRZU33x/Y3uwa35rPA7GI50gCgTh6Q9K9+r8uM5IfWOjjKp
0VU2xEQVkPgjkBbkStBiGE3o9LLB1RRo7HWw7iylAtVxYNpQcjBdqPiwdkzFjp9m
TML1OBiJwrMZ/oQ/ZVxxwSV1effpbdo9rNEwNRAcDuajIdc6jxdx+IsNdc6RBpVt
Y6oKCzQJoC4my3rThZQnhP58KLcd5y8L2OQlJOV31pqc9r3qFaokbqufZ78xwRog
gDniFdWRyiQLBWVWV/B7xsR/3gh3AKvH0w2FLpLjUpuGp8OE37/n22j1Vn2zSX6w
ugm6ADOYnbtAtzr1oGQ4e2tWR4Bq6egnAIr9W6SU2mPcJ7DspkXYUMNzpMSagDFN
LfaV3TQn1rwchQoOQHLrq4NqrQGVY+jSOfC9GCs1ZSX82JIkcL1AeWGsB0PIeFPv
TfFArdhpOI7ZXnr+QD2DsUfbEyLwvvmhgykWUvRW+82JIZpVzXQPMs/fYX+fcCVw
u3mUb0m55lUi9KhmNbqDv+Tb0wkf4G6Aj9vmBXK+5f1CPqpbMcVLk8b7Z9M6yDX2
cjnk+1sZMYANaAEMFdJenba9DDQJvKF3ZbOOv2hCEk8UlRt3R1yFEN/+Z6qLoLuj
cNz1nqvRNfK9JCMwuRz6da0UwSNWBiSLAQdzPExPCq6BeT/iq9TlyGY0Ct7TAp0u
axIJoQxnOuddHhNzzO9He0lJUAyuMJ5dPSyUeK+risvP2phq65KDUbFZAQr5EDiq
F7SVw2GqyjFX6yv97AiWof4+3DzaraSN1LtYcNQpEhklq37bzLvZtcKZsN8/XSp4
LRXPraqTfBhSxmkPNdYqcW5k1nfiwp+kqBw7TNEYE+KEF8TUMkJjAc8xO2/rWb6C
gjk/l2ra82vP6VbdRKbxeS2oWGFRuBDm5ZwZsjKN0nCk2Bi2LfwEH46pIvmXwmv+
IaBANrMZ2syC1vdhU4HOfrCWWCe5k3bviVg71sg3jeH6QSdcS7q7lE7+1LNmOyz8
vhmJdDKjA/vwLs5KbaFuO3r0Zak8IrN8DcKxHF6vwcNrrLVmTgNLTwQ4Wm6wr8U9
5Un1h3DTJurtA8M9JovJiQPQFVa55LTGMVh8XB9o9wQsCi3ni0JI/v1uA1NEvFRk
wrJJzdIAPSfI9usCavqEBe7FAkiUtF0kjiXo7hxNpqTsIqdyPnm62jMuFiwTRo7G
4k7Sa/SBCBnx2CDcCSWTEybUe/RfXIv1RMu6DEuZMVa3PhI3rM/ux7K1jDaDJCOB
JOeV9d7ElfKjMpriTE4eqXa+DYtwGaV77d5eC4CKT0sdUaqVE2tZPqCwU5+67Qig
NxfZuNPtHYVeSRg+dS30goPkC8il4kmpioiYZvVdwsOuz3FX0pA+61efZnMzhtEi
wsuD5srw4V42DnQEQY0a7WInGyiFd3z7zwOHKAwXSKHHcyOxNrFqXBu0+5tZugOc
qWQCp5U7vcWNJ1qyAvSXOnWVQ7Gzlky2MXiUEr5+eZTW8N9ep3vW3cLgbAEHb06w
YpcQ3yOUECRpXPjVuDV0nrCDXKCGrRtZyw6sxuMZKx103Jyx8MwsxEHyoopcm46v
BLCJEk630zlx3vhER/GDC6cKJ1hGZTwgddDxSp22RCUrTRAJNAZcSStb1KBPt3q2
G8pqSsaUuovq56wp5u/IBek+aaSLhCuIoSJT2f1xEXUC7UWxFhMdVx+Lydw00FY9
Smlw7m/lbygxI97YKv4m18CzStdajwlC+yccbigQ4lLm3p/tliekY86NhT6tLaAS
4OtsKapaoAun/hySnoCpOwzzbM4mIb6UkaKHy3eYLKduYgs+pdotjw9XKGMx4A5s
wK0fjjojkYnJPuJilXIBAkoJZlA2VlEp0v9+nlC/f0BzXQRHsZdkCd51GAjpmCtO
7qRsUMvscvQguMKX4Szdsn3XQ8MJ39yu3Lte0s16KLRyMSBgnsdt027UBmlezlqR
yHMj0liQPHOu3su42ZP9/HLzzhiS5T5KOXWds++RLnvrCtW9mvNj1FVsVxAyOmyh
kggV9l459+w6a+TJCKKBFDiY/Tv7Nyq9rC8erpIlAgBDYJoQMJsiSbGUJouESzNs
tdxcNmIZ6HuvEUbnTacJ0FD6w1vVRtimH4ioEKcpum4+1iious9eSbq9jMR3QIG+
DNBbp8qeJLxpDzBznN/ghWijRmWq9g599D3iE58yCZ6nA1rBLoBmfK5EtGot8rBK
6MdiWYAUiIcS8NmOHGZmILpynI7ThBxhnkzJs2RKmyBmep6EboNDyFl3F59g1uln
+VXDyZkab4Mqy9xdno4qt0vuu23mm8+z95pqQAUiRIE53YiXylXRkuR9egq7keMS
4RQiozVbg5LyiztR5SdyXX74pLv8Z9P4s4RHU17AdbD0DeyhunpgeHU46ME6U9YR
Zm0rrDURofBGu10X9649ziwNp0MMJi44+Lxb/O2UnhOu8M/MIs8E86jWDSPIaSDm
v+PG9484x+RkBYXnQksbB35iu6Z2DJwrds6TMom3N4fVh9lJ6/S4J6sIh2QLbdUA
VpCzCasUkEaYKj564TuCTA2xKoPBpEjN8cmr2DTOafIiq90d40hxl92H5aIp/uEA
KRRCwBAeSByALg02s91nxBaz9X0xQ7VvgdsZONyt+jAfmMn5145Hm4bKnYtSOESZ
3b/SuAzI4ChoeqGssGGB9s1ENM/xseOYdnPQkZFwTOct8AJBW19QV2EA2cred4dL
/27uOQXBmTMq1nog7+dMrFZUhnPrwdhlZmk5XanH96RP6eRPmWk4zlTU9ttu11JB
TzKO1kGK0idT7ahRVwBo9/HG5+ntCXKLSsMpDw0Pgsu9O1bXQ7S22uMEpjf1/I90
sRukfJ6zm7YP9oUNmSFxMXXV9WWQ3K0Ikq4hJvL3ybfHDn7PSexbKCQ9PqNptxtk
z0AiKFmsv0gzQ03zVhp4AREpcY82P9wSs3jhDWVZ0Bwy4wcYonw1td/0bMat69hr
tiAs6G11ayNUPthVKpAZZI9qXBPy+Qi/8SwhjY2rDBKT9GBZp2K/OmDtKR/tgR6t
PMyq/9MypioAnf4G0Ux5WSdNT0Ly3KV8KzdW5IlMC8vYY0KatcgyY2pRibCn/Cly
ZLF1pKG08clcIh8WUsRBhCvZO2nx/rxt5ikcpMbqOVcQ/DncDQ5o0nJRJXB87x6Y
O5t2p8hAOMDyQM6KcXGROI1HJb+siCEjR8zkjs7rrL9EYUq8GXPDPxp6VYSqwmRH
jhTqRoGDehBBU9t036LR8oOthWISB/a9KmqYCLrRNTzvgHpicoxsiFe04uPLO3gC
WYjC/OJMcYu5czXiZy4FWiPjb9P6GxfwpJitRsURiBe+IILusIz24lV86yZSdGdS
3HLuTmyT13fVhAEkf7ieIfZYCnBj8erh5rs3keBpeKCJxQy8dHh7aJeH/R9YqvGb
eW/X/O8T4OauY1y92QKLrE6M2lOGoQqpyO4Kp/3wUh8JpVsArjhrQG1UMjbN8sHA
3t5et2utkVdMZdtAQHRSf1FmN8YYlKKCQwxzOkBO5DX2/XsFzD+D39pgYj6Yewug
HV4EuyuxVqzkTv7FVdDn1orAJicbJ6WFfPGfXXHLTvZ0umP4dZsNevtkzDdMHK7y
MEe/zURadHKy4Y9Z+nwd6565DaDUWaoxXtzAjUYjCVNHUCOKt2DZ2QKhOtqYchro
gb7X0ISdQPzKvgqRbt4FQ9J6Do+iCrHwMYW4/WASzsGSXU4bVS1RwtYwhRLYCjrA
AsW1T1AvxG4GSAZcA9aneFp1PMF5boy7+ezg6Qw4zojFpi6VNLF+PLsxCK0hBJZw
gZeMFyN0zCfTMRSjg/79F23pK9LJOs+cDcLAJrN7Pyl7kCzpltV4umE61r8baIe2
uGdUOSog5Hjx6JMba/yTEm5OULA3DAqd/JA+YT98Z5ENnOVS9RcQcimvD/yoa3xa
nHN+j0zK27r6CSJKsyW/T31LHYQ+Akq1IEz/d6RPNFU5n13GFb5lxOQWNTfRibXa
8jkTFk9O/OFkHCucTX/JBuaU9yUZToksbgncFcBALqXiLaRKRoCFxmRmfiJH4C5q
yhCUOAWI28eHqs9NdN696MQzplcjz4stpjpjbsOGqmcrfaazNb8sUzZ9fiEW97eV
k1gSYKu1Ur/h7vkdQszon3g0R9DiBb6hPRSj3KuCdIqXQ0NSyUYKR3j4oxa2HJUO
4obzoMYCWg3tPk0KcSNzj6xinRUV+qo0+6HrlO/LKL1SVSFeVTyRfqIKf46ak6se
nMYcdw4Ovxhw9ii0IHgJ5HBFuU2Ejq7X1nCg0kOo3Xk9/zidNnq44CfDtn85gONy
+oRY9D6lhRvDSdXqCPgKII1rfgLeZYnrf/nyQ87R+idJIUuEpq+NVFoaIprH9/G8
4st4UDyS9jiST/dtwFEM3ynI9N5kj1zzKPzqaA5oQSF9CNJQ/ax+RKx1mKJturYX
XMA6TVG8mNZ5Rvc9R9p53cygDkzT88LZ6DGYG6GoAbGoPpkr9jfQh7FMGUI/kSxZ
KyKRFP2NLl2/tMo6td3pfber6Yat2p4gSBdv5WzZ7glH2Xyvv0IsOGjQBGQKKeLJ
NDiGyi8mC+1oVHTu/AxwcTBdDuBh1M1Xcxnh9TUAGeJg455oBsnVyUdNRloF4CmN
iSpIjcZjr0D3R4s38wPKPYxp7tFErWRWbJPwPjV3Agrg94bSeqrHrUGtzGdehCm0
B2InJnInuePRkFydV6kOVxtSG85wtrOoe1LIGWBQ2ec/nSr1PM1Wt8vLxLtqAKDQ
s9+QD7CY54gU6rHgVm4Gx0w+fi1VDpcJvjOk0BfV8FxXQjJZxA3sZ4RBM36XBSaF
BZfeMjmao+kTaswwK+GRSIV9zt38dJbriNmoaFUlk3gxzbSEla998xTRxTyHAGNf
ELYNXsj8Ps4gwKnoq2nFdv75UAV0Pk0WATcytWiM96OAEsk33KqFyT5VB8z24uA9
fZcFYpmCJpVt8q0v7q7Qolz17Ni4zGIrD2t/15oXSrX1EhIGeY6VoIkTMkvC4SnG
oBLeYqAygo8TFmzmha5gcU/6sag+vdfcurH6zFfKOS7yPlYdkpkmwZHxUjO7LU8Q
GSV3lGsYJRLTfh0J0CXw+y9UI6uZ4KLKlcMWi1km+VRqS3psnZWV3yrvI6TyY1rk
ptZNxrMW/1rEXITWUQqwRhw3eASaJ5ZEb3vYv43VM+wXO3j1K8HqbdOXQjKMV0EF
FuBlp32B1lRtWdqecBnCgkIck7NB04p8LoLn+GDCv71cNzEbkiYk+LiXRyOiI669
vH4UcDTv+igxp7rl2bDDctYu+zDtpbhvMeRsEoUr9Wsdt39X+qAFNssVBs1qczPf
NnZx/Vl3eKAXAL0aBIC2Dd1x7LXP7eycg7oHB1UwgzIvrwEiqnJXW4wDHmimjPiV
PL+/iB8pMQYT1H+Dud7LaJQDRnDOQjCtPWuDMWP3NnjfFqLdViPcEaKxRjKisU/D
dukDanae93VvqSk2qW/sDLPsEn18Eku0MRCTS4jZbQL/sRp3QtHWbHNWvKWq6S8D
/UcerKRY1kBT4kZkdbCyudYIuQS3DlKYGro2MD1YuiYPht8JrkMvQRaiUtsi8ohk
EKUDqkSSOdnC/t56CaYEvgHuSVrLOOI0uC3m2WScp+JIHJ0oyJ/8pGyqyhZCbQZA
wR71cTxVHVEv645+c/3BA4VW7WMNGqO7r4HOtY4vQskovF10YlVK1IUdg2s8lYW/
p8mG/a4lgQ2lv4uvZpXziUyBVrw9ZOB/u7AXwqCLhYf2AB9x4urm4QRvcG8+O3Vq
NhWQIwAfPa6ppTqxE1jP8nsIdoRegaJF7kTr7qUCQn7YAgxrCplgFMXb39TaNmg9
mrdAaaLzMxXk6i5iyfJbOghSSdsDyMn5/CgZNxm4U4GEx8hawcVzQPT70dCA2RVp
0mZNSumQGcrsS/T9VDKd7dDz2u7w9otEIUdA/3N2O5u192/uDgYTnMCiClfBEMtA
8bKHRAMPjzbpGPXDlNfR2akdyHWgLHsOGuYejs/vVx990phRYSuXsXmodqlnEC49
6IToBHRadqacRtsdB+/VIybQQvDf18GmePOyltqi4fr06dOTx1ZYRDqgxybFR4Az
hXCOBdwbw5b5nse3smauHE/LtgdYj2eJQJq1Cgb1wgqwRyWMXiMrSOGjzn4jNw7k
KJGuZ34wcN+Q/IwNNywfsyelyxbE2BNV9g2Xwq3vPmYA/oD3Zo+cAJVbhn8GEyGf
2AjaCFjOVZebpm4s7BnsJIjBbzmFVPqYj4u/8Mmn7QlaVI94Xw6M5LkLSpKChoRB
u2uVxlq4lQrlmLjOhs92vH638Dh2bwf8zqoLdsqscRHv/ClZK3Nd5z9vForl/oE7
xJIYrb8BhewRdN89Fv9jfnCH07+qK4VeZxy19VXhnEP6eiCg1rstxtFGijUCenig
ZXcYgpQIXSBfF5t1JSQwrDjBhG/dEXxB9QHF+5MBlUF79P9qi6Gup5aNz3rcfO2j
dfyRB3ks6/RNvVv8g58OGVOL/Qb2tjGfSF07WNDRi0gHb44nZ8U4ujPul80IOjgc
viYdCwRDOcE5mTcgjOjaw6Mct9ojwa6XaoDqf8X+TbGmWkB7ei4t1LFavDznlo6I
r+qobO+CRWjEjIUTQFKfAHv2fq/w4Ja3pYSMpEW3A/Z0559fhhGnJYHhwCCBWWa7
2PKDnRZ0d926S0BHoAOrclc9yXgdRTmVWW6rF/sKQhuy6QUqy0R4r+Rx0J3BmqRk
CMmTiyKNr67jX4mkuae2gZLG/1xVFkKlFdb5RMPmAMptSO81LvJI23a+40zUWIwP
aY3M7CaBd0Ef3QJK3L7MM+WR+1Yp7MluY3JkX/q5nWUAFX2UO2F6UbW/UmtUREPx
UkNfpnS2wXUdmkFK1tW9J99HrENc4o7cHP4D1mmn5YnAbK8ruNSzvP+NAouD4bze
fn0DT7AhNdxkPDRblXacEva66msTCHtLURHFrLInsAgAeI4t7VNqbn5gJoWAn3q0
sfo5Kivd59ZiCuEq77nTvbNgge5NJnEWA/FEtN5yaZeW/X5qeYC18jqTj8wrwlp9
bPNG0FgEoShF5bv4pB5mjIbGWOwFpkKgunEzkR4BnqNw0GdViYpjH5IDC8TNUxqn
LGKFFELrXLhetFTxztHPNH+aYhnzKUNDtvzAlJVx/qrlqq3pDOgeyDTegSG+teD4
q7yDyHQYvGoz1me1a5HOomhSLqaLYUVb9k1EOtHspJaHIVfC0RGR7Ig/qwea+cyR
t9mb1Xivbr3od1rRmm+fVrcfIct66zmeHmR0UL94RnbT6+OI9/gYQemBpTc0ZeX3
ULx1yV86EISRbbq1uISLoObY70VVhkuJlvGgpj3GmEh05V7LB/EbGmD5PUOV6mAo
pS5yY6nVWx3NxJmXD3CEaaQbdHZCJ/rLmZeZLuoQVRBRXDrBu7NYRWFI5KQU/LEE
3vJNRKF1Td/Yl5oA3un9fZlpGImHfu+snVeu2/1TUtnyIUT17UAL74Plb8RUM4X/
gsQTqBvSy5FpaZCWXU1cQoWq2+pF5aJb1GHRp8GNExRLMWPxW9SIxSQzopDSJHdl
RtuEtoAIiSJhmbPA4HPw29+Dh388WuKFckmMDOiTZldSsp6gVYBOKatPOihSM8a1
1diHJEY7JGGjSN6HSovhHQ2xNK3R8ylVXAdpqGHHP/xfeLA9OH6Y/ihxGG4cwZX9
0UYDwJTfg0R4/0Rlw3wi8r/qlUq4Z/mS8yQj96gQ7Wq9UnVPQDA8s92jMDQKzGEK
EAPMe+JpN1hQEffYKB/rjoKc59dDi9ecjOJ+IBM2LJ7lBCOy44XeG8n2mt6egrXw
lQY9sVyphb/Rw4T1sjCN3Ly3T6qeiqLVy1sz30XOvsRVLPsojE1H+pdIXny9QSoI
LDBQxitaEAqAhqjePTBuOF6oZzRkGNYkQnN/hAYvLTV77kTY1a3EJvzFoBgE60e2
yAg73MZcLcMh3FevIufLTvJ8RWsE/w85qUFez3Luf2LsE4kiyGP+McAyvKdMFCTQ
Um0dprb8cWNjp/B1pXq8ZN47vyyLxmPrAGucGl4XBtGbDceT4I/UjnU06YBxnBCl
1HPL6b2Oetu2F47gNSz621hOO9OKkNbcHKJQFqPH62qGmrW/XF7R+1AkaTctJKb1
aJdQGJz1V2xxWfN7bidjqAN0srI4M0TzpZcF2ceDOe+ihy+uogF1Jsvio2PHrRAl
MR1+viEOI6CFQtAh4UIjB7cdzjCOGOJvRvnfmvqU+GV1J4XkI57KaQVQff75wnbW
7KbVoP/4kCxGekMm7UHw4K5JCk8GL6oxDtQHplH6/nxumrkzpECziZMRnYnLZPL4
/8Jn6qTvxHGENI5F1NicRh2uVUFYUZnCwzqkVUP0YdpmbhXxnujACAMp0fgIdZxJ
D+irRp42GcSbDLGhyAOxoQ46CEEGewBbM6jxmWAfsoSDC8ltS1BHVfJgnj9JabTs
ylMpfF5cGYy84t7wtlooEVT+8ZiFGF1XPwKu2NjJCURQymRcF/orQEIDKOIWjj7x
ji2TjnbccQBs39XkVPzCzBEmOoQDUlG3vbrIIOn9U43CaBw6BmROlHKQ5sUMvlDk
ofzL9EYdU5qU7pGlm1/Bjtarv7/uJt0m5L5RE/Hkvio09N6z3o6JHkRuvRHPNWfV
iQh2qbD+oaEY4bvZDDecsJ5VyA/QxDMqaxfR3H8eUGXBovHB1JUgQbHR2WJi7Age
DuT/62BtKaFciBYZ8OjD3KikYDqucv3r0/dT6pdHPPlZyivk9J4WNJY1OQAZvTCu
VAgt7cKrBlIlvpHSv2uf4Y77uLQouFB0KH7WH+PAcj9Nt2rO0RxZ2YiHWn8LpViY
QF+uqYx1xxjk70AFlO4bMkPvDlcW9WR/JkLdUXO61cwl0UAbQsCCh6DRYW6yBdHS
FZmPOTJa/ra3tdzhX5UDgCK7l7tG5Nu7iEdtiFloyK8LTw9XXH3hJ33HhueXURE7
uLEcoLyWDK9PzZFcTjCCEOC57Sijbcf4nDK0ewvDGfvaExCcVmpOebiddc6BphsT
SO7FwYv9kGWfd2X9S4vw9G4VreYjSJtAQO8kIEjuwYcXxsfab9Cfzxa1tpnRVlT7
gTbfq2ZPyUCq2TAHWURzEqOIZp/EJzDcZOD+VwBXOS0Mc9K6pHGcTqF+fqllCFjr
yorXcFpc53GJndrS5xD5Qd0NHZxkkaTVR35/0n0hzUkxPNnMYQxmRYJ4IGlRBv05
dG1FaKV0felDtYKcAleZmIlsEu+GlsVnHUo7QO8JteHYPq3v22/g+9lLauGLJrzO
KXfpY1F9gOqgspWtZI3pjsyv9vwGG0i6Zg9lAEJS1iN1Kk6WYl7yCsoQgm1S2kl2
auHAYNeJcSW1kpagArT5X2IawU1drj+yS8n16c9hx195+jBtHO178hK3jFNawgsR
WVtUT49dyxuQ/NBbzf7Uq+D1Nz5HEGpTqCTc5ZPH8mhzNWAELbT0vkBhIXcdzsmH
a6HCFjIgfI3yQDfPBHf7FPGOXqyiRyCspzcP0Q5A4TFVrfmTmtwoQsDBONT9eT6+
Bcco7/qYXCrAVVAOYrDXesi5fyK0JxYtZISJJWxzZ8ZzMLMi0P+jj5ME1Cmq3G/F
Rxr9PLG3e6k0uSS5MhZApCfcOIes8zJEPVoSsXRBpv+qdaNoUX821AraeDziTPMz
yBungXqsK1c18sz6ApLdP/vml5pKOYFNE3xzogtktltOjYnq3jdyLrjnMg5utIO4
QUNvniED2e7yEBdjbNxWGa3VWLOoNsUb9M9O/P5bvezBiEjioZHeSxwYmI7s+uW0
IHZ7aI8nwV3/cxY+1/keV6f2mUA+ADMGD63XplxIkUvO6LL+3dF8jKe/Ta1RvlCe
rxJTyZUKZOAryKJvZzcpfNHmWg34TSDLGPwiLgQtkGs39VO/8wuzuUuFuuI5mlGC
8mK9L96JfAEOhT3OzBHXACuzYSLQztrraHY5HvTcumLhKFPhNBmNk0XYLbCifZQz
/os7JMF+H0ucQZiBn0GVm4lfWQZhe9VFojmULoHsY6xGVvlr25zBqd4huJYY6/ou
JLlll4SvPhIAtfGu5SiWR0AXQ+QVVjeyhVC+1Mu1d5e0Kz+Q9g6ZUb6ByOP0fHkD
1/RH1jKeHdOt9pzTiFN5WBEyRiBLINmISjk+cZLVBeNiolgfmeki+2ATADTIZYCt
35CoCWyX0XmvKoMPJlGpgKvcGSXBv4Sc4XIeNV8YGrVqJ/wI1xsq1alLWCPRNCB6
+BfFuExT800pNcpjT5w3Gt4y+d+9FXBkLl7Ofvqsu0q58JJIjJ1+L6ON3G+yXGPK
TzrBsnNM7ZJwqtAcniMPKf/w+zxSaY/IZsLUeX0DCu8PNdg0oqbaVQ1OSc4NI1qT
kbyMgF2c81LR6ePfT1zu3o+ICwa/DyWoX1hBERS6f83qJxZWOXajGGxCdSqZxukw
zftD2a3w7ulaFWUDMt33DFpyfWrttpoiPifG8Ho+1/IwJGBl8iMRBmurO48S8YxL
oLPNNf/8q7b+64/0gg5xaSikCxKM2pG7dJx8elvqRhwRKu4Gg54LsHfXcMW1RzZ9
dLoNN6JNMnITs08RUCaBMiMVspujTFDmv+FAQBcZvKBwzpTTfPFKDfVcdpDMcCrG
kR9KReFdgYOVtXRS54UH+8TTKz1DBngwyfuakwjyDV75R6vSzLOzQRN6Xm714cM8
EChbcebHKSkUKa/z7Y04YDibERhAB0QP76gne+DnfF0b+XiHIGfI4SU0lXRuW31b
dcdhIfD4XJC5q+uoU36+xnJ6The0QI0eTjM98N7dl4WAFelzNNW7GK6xhqyoEEYw
DOEa5A1yx/jJMTh9twp+dWmP897AYLAm4fwtP8OXoqZDiEx2+XC//T95NEGKDF0R
Rg5VdiuQDyjaJFWtEQ2iYJQPeOjKCuOakNOeyz04YZfLv9QX4tvSU3Fw4oWZjBk3
QJ2+JNgttuFi0/rn6QNFIHW/2bK427qJ9zTzw5rm1d+u7DQmK6GGopeNKd5KQda1
IWvOpWhgold/E1HEzcjcwim/2O91USjj+IQYA0LaNj8AdnRg14HMP+Z3HYGUXerO
f1L1Dg+sPeJY5Uq+/mtgHtW62+6umDNoqHbY2yHbZTRPnM3e9JPilHvhxsyjyPe/
8OhBWtVwl5EKzsRAD5wQL+O4gqtkZGRQRih/wjcyrEGxzd11FiNWIp72LTIp3nkA
Avbv+7VyZBxbLfDVWFDepTbiSpnSY0brTS8OJImHqFnieBFtqcy19N+FB30iTW70
iSk7eYt8GLZyYXOmdnSO+0F1o9GcqO/yre5mUhodmWkw24bEBh9RTx+bigEJHisY
GfILSduMB1wHeqmNIFH0if9512tlA3dOxPj7tW/Sor8vRdAIllyn5ikcC7b7gDVn
I3hprU6VMoI6Nxf/+fYBJSjqdBehprc+EqjcnC7/H773A5HKyoUK+gpvP2wKjPHF
5Svefq6yzfvnaZX1nl6GJaP7PVcHeoBWfwooxaOzRK2+qQVmt72jaNsvzN9spiJp
NM0WBWppehxk3iEIr2QOaXzc4N1dC9uBuc5zUlHr+7GreAjmKndGqS5bBRihsqvb
aNsAZV8KTtHte2AnGRNoUlJDwF6ltbSN12jZLYgZmLadwm7s0stMyVGSmYeelwkC
RgAapolAdsR/ylyn8rOwqVZ4tjA9FAF0RGbsQIvWhAFc44W0DJ6jv/d20XeSX3jd
7dmth2z9UwG4K4sswqUuZu5B7T9mdUFDctHcK917LUzMP29i38TYz9sYLllkY/3B
znNu5x2H6sjyrn0CCy2tMoei6iqopt52OM/mJUEJeQIOulb0XWzVya2l1AFFW+u8
30q6Cz8rQ3AtnRdFHmbhw0PK5Msp9lw+DVxsgo6TSrqm6h5cauxp9wFIha7me7uq
yiUt9KUgjEA4AuBZbYjRcyY2mW3lY4KTJQejYAoBoq8ipg7LbICj4mhaFrQD2TrR
G4FpNVnPnOCqdO5H56UXMicGF8RQrk73RAGBGfMozN0m5dooryI126cqGeeBg5jP
WRm5ELbU/gkbz84eWJsykkyl6HSklecdTknNnt09JpVaBRiRXOqCbk5HarYfvelX
x0DLKPjiBxUpT3pjaAxLtQ2sjEPnAKV0IXzxGHgIjzJXaehL2zhdecoY6UPuYQVx
DZT+3afvWo7DYx5IIVsAad2QfYngz2kBs011EzSMh/lOlSMvIeMybeh6MJ8d3D/l
DCRi/A9dxjQcdrWGa7GG28tClzOLTqgOG0so17NFAAhxaRAHF+UouLkU5yaMRMz+
wCk6h5RO2+VxSBr7W9uChQMYTnS99cAT4QKQJnI1JQOewa3CEnzh71+YtuCO3JwH
7/FZUzbziMWNLZjzAyAwpAoEc404vRVA/xXgLSMfhmMiGGKT5cKIrDlVzlvpjb0p
g+jG+0Q8GrtdmjYj/JGXO6sw5GZu7rm37brPtfZb3doBBty1a3bEH0DQNtJetuEF
RlObtX3PjzIPxgK4D1hs8KPA1YrEiEW0O+jLcufIsHWnBJtqSk4DCiD2lLzUzIb8
aIpzntavjLEst4NSb/t7Isi7hSIQjwaN8SYtpOfQI/XqqvdwmWcjmOCtCUMR7Xy6
9BJ3gfHtJS+dlbyNbwQ6/maFrul6698nCcOrwfFyd8VOLvqNVcMoQ9TotqPa7bQI
5lO+Qn9yvC5Jq0R1swTtWlbGuHlBArfjyk/VHO2vUKAHQirjuy9rqVm2DeHafZ6v
+X1Oo4i0EOJNtFnU0C8HH13Nn84cXg8K4TXXfso88F4KQvdMUo7mdqPDwzrJYBM2
Jv4Kf9qwOw544Bjpm01W/SbFSY6b/gzY1xDUBhy2ogNpj17oS6hZHeMAebUlDqLd
lF8zBbcOWQ07Rus7v1r27ElPQ8ADZhx/KsYF05vuWV+EmSjXgNieQ9d34DMrjoO1
napTH8fAUJIjinLQ4MpUtOxQ+q4+WUMcA8sGDC63Eng0taWP0sIkLfmI5uBsG1bX
WQWGlaQ1FSmiwBf5FFNpHzENWPvYm5fKofyEN8XUa1JnZJzwsiYCGed0wsMGfcpV
tmhHH9wySUgqAZ3OSJf0KBNNHYiztAlkB5UuGjeL1pH/9uEKRSdL6KUZtMHqgi4b
H1pIWuBEJfCldUkZWWjMr5QEzLxB47ldi7gwUjuMhKv2Wp4h0xdH9nUeo2TTRs9h
h2zClgiN7pm6X/lXqiwiVn40wMmVCu0oS1HefMryT9Mz8ZHcN2HW3p745KPQRMtE
gPjDO1w/39rXSySzg3TWSARW2yVyRkvcASHJvo2o2AYZMXDvkmSUnOLvsZTtILEc
RSvZOGhq7ZF4m+U9fGX07ay+ilk92USN9I2KH7vLIvmFFh+wXhdO3lw+6rBI9Pky
0wxDxnNP44YLc94uHf0moBr/laL7jxALpCj8rMPGc+7atg3Qh8R4AWPYoK09b1tS
g5ihkO2uUjGxHXPlIL51YMfOSZk+5qHDcft5c1HCY9U/ycjybA6isdEj9I9LKvDP
T51JRoqXwJG7NFB5Kcp/cXPFDcN69HO5XjjA5t+0zaQGEvPi1Susgo1ssPT9GKBB
e8vBXsI9NOpQYGSAE9Z+NCwKB+tnh+pHdfY/b+DJIyYUl/ChJ7Raz2MxnmrQ74T1
wSliNHjZiAczxVPxFvBplA==
`pragma protect end_protected
