��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:�1A��"iOWV��=�}k/�+y(�&5����e��b��Ѵ���$��З6Mv�Q�Ɠ%��oI@�n�gӧ��������P�m�;7z��md4�>�/�-{	z�C\c���������R��X��bm9�M��HW��Ϫ��s:;�\�2���XY�3�h�8}�������e�5��^P��֜� >X)��TN�ѓ�@��!��T|h�����0C��-L����?3ua�(h�%h,���1�(�=���TnŪ��;�� I��f�2�If>h�H�NU��q?ޅ�wud�`p�8���ۖ�� �I��4٤ EW�
�1������S�?�q1�&"<���sk�*��TǫoP�JMw��U��|��'�u��q��/��Ć;�Y��/u&V�O7��e��Nc���&D`�R;�^]�J���E��
�^�����[���U��W� �<�ۈo����QB;�j�j���I0���JM
P�5��P7\풞�l����w=s���<KQ1d`�\�"%<���4��o�G������#�������tg����;5z���M�R3���l�(
`�;����������"t�;$�U��b]]/ˊN��3�K�I�ƛ8Byso���__[�אּ��O���đ$,��b��� Q���j���3�&
���
*�>&T�����2�o�q����Bc*�-��-j�Qd�]���f��	��?�N��:>9i�L��a[���ml�o�D�� �3�ݜ�cO���n~	��o_�b��ɠ�V˜�c�o���Zx�8d�<�KS�p"��1c��Vd���D#B�>18��:�.�(��3,i�ۺ�qQk�BBp��J�����Ņ���v~�C!/�~۵jϟ�ǯa@��7Ö��A�>jύY���c�M�R�M����x�
��t9�G���\,�)DE�i`�yc�,{��n���no�I{��pa8Z. ��#T��MO PH�����H͜�VEC�\+FQ"���C�ajsO1a�9�t��Q�u��s�mѲ�S����H���4� �X\h��P�?���:E$�x��_,�U�y��_%a��\�ӎ�ߺ�+���:��}������jKj]嚏ߓ+����5Pt�흟~6���]����+��&�Y����>��O2���D#�,�@2�z���y2�Hsl�%G���,�PGF��JZ���'������(�����}�G�b��xX�d��>1_@��;-��l#��VǒoGn�F �a���yz�d,���3�V^��s����#�p��[�<#�#�V�ra��&��!ʦ��暄�,#���j8ܟ~k5Wӵ��: E�E8�8ň���Q�b��:�9T��	kZ0fC��a�:���.���Һ�:p3�ɑ�rL'M}�͌dGh?��
.X(k�_eL��7��Թ�~��K�ph�x1�m'NC��^t֖�c���q�=���>�V�eʖ�0�n��?(]@�IH�C� �ΐ/�Xf����N�[o�k���3-dpw��V @�̥rV�T���צ��^��1's��)�*b���}��~�l�ۓ��Մ%?As<�4�<�)1� VOVݚ��SY^��B�7�x�Z�����B�>^�h���ֆ���|���x>y�nA�]ɂv��b��݊Pk���,*�)V�v�k8YQu�2R�7�e�7r����/�Ӏ��`ڎd����$؟e@��R��ۿ5K�=ƽqP��{��i��N��g�(V��Y &��CPFG��/c�Q��:SN�.�o���o"�JD�.R	?_6��>vgjb� ��/�d��{k�.G�&37��y��o��/v�O_K��d�ܖ�����%�6�Bj������1���ԉ�|�ZS�͂ʏo2�y>��׶�t�ԧv��B�m�u�A�%ӎ��-LƃC�B��4�7���4��#!�3\ sų�z>B��.�JH3rkE��#CrY�֮��[��u���
�2߾��� 8��(�(@>Ĉ �ˎ���$|:����=�
��J��`a��0��_ݬ��Y��tp�$^�(���/SZ���dvF�3V������M3]�lL��m�����g����G'�ݛ��e��L�JʐO.���G�ɂ�Ơ'��ƞ� 	��W:;�C���']0��¯����_�b��Y$W��m�\HB/,���N�C����: �_稕�0oJv����"��� ��X���ۻ>��Os>i��J�}k�)=�q0��2��WE$�`�H\�_���2��pm$a��[f�X��S���<%���#ʇ���vh=,�,F���@�,_	{�p$�<"��W�
�i�������`�� O�#+Zv`�V���ԕ�* �a������	�)`��/fR9����՚{���u!Ƞ��c��KM'�����8r i<lC;�{�X.	������v㠺�#A�5��@��2̵��޷��ͽL>�MC9V��M��Ӫ��
�10��u�T�:f-s�zyqK(]<pI0Eݽ]G��+�48���Yd菝����R��i�Ԃt�vn���+���U]�Mx�|�?�����~��b��(����u˒H�	a���+Cv!S,��k��K�d]"�2�`�1�U�偀LOșG�`MI(�Y�3F��κ���%r��l�s?M[���-��"�X�_4��m�;&&�N+���Y%��LOx��t��f�d�	��o��`ҟ=zY@,��&^��� �*�6���+~�OǦݜ�V�A]>?ȸ�����(	�w e7��貱��k�P���ܣ(���rs˔8?�X	A0�I,�����q]\�Bv�gO�R߇�.��Rw�`_i�'#r{�^��w&��M��2=�����]9W;��G��r_�m���t*+�[��̦�Gvv/��<���%S�d���W����$�	o�:�A�G}���;�����.��[���6��`�BU��%��VW�J2���G7(Mƍ�>�4�f�����3#ѳCfG�s\K�v����x�k�~����0y��{"�����ꕥ[�YF��ϰ21"t���'�yz!5A��/"�_t#I\_��.���!V�F�V"��>8W��+�.�aZ[r�~s'l�t���t	��.4�j�l���u-��A=�iuO�3�$uv+��sU����"�~[_"۸��C2^������tG�#7��X.t�)�;oƶ�0k"	�������ã���l�Co��;T�v���pG�ޓ$3ͺA1�R���n�g@���1�Fqu�z�@[D�^��7]�J�W#%�)޸!��xWӾ�]/��iS74$k[9(��`�Q%��pX�i�(���Y�;���T?f�c�l\���+�,=����k�qrM�F洎��*dx��� ;�5P�ͽ�G�ԩw8hЗ��{���I�!	��5!�qŇ�u%���w8kk�ɅpxYF�m��nL�%�){�v�Q�r*H�����F�,2�R��F�,_B��l�}��Rx���Zz�UKs�R5�9�ңpK�n�;�E�8��s�"��v~���{�y%�4)MZ3����T�twM:�"ݮ��^�U��۔���se{�rwY��C�ub���5n����	޸�Hr��% 8�ې�x���I�Y?]!����A�,�,2Z�5mT�q�����K�@F�F=������W�IE�a���川��ݭ;i�㶤���.j��S�����֥сrj�����P�f���bs*�������aɿ�;Y� ��z�W$�e3��h/��
�v[9�c8þ.����.!�KV
���d٠-�V}I��v���0E�h�\JSj^��6��_���m0���h4����9?�>Nwi�������ls���b(j�mLZ��ĵ���zs5w�	]f�̣�|D'V��5FF��Tސ�x���k�oz�����n��Ԡ�0X� ���|N����sa6Q�LwR���e���AS��&�52Ƹ�}��A��=#;�d3��	f�p��h�	$�����ыR�:�\�_#1�	W;�j�T㥯��ijx��`�C��&�dEǿ*IV��1��4�� ˮ�+h�v3��<d'�}�M�'�R�#�)���MA̞Q�n�ـx�X��h���t-��Br�.���#��̻���п�z���Ý����@q�}#^�ʍ��(�-`���W��O�2��u�1�=�b"�<������o��\*�3 ��렱J<E*9��гNRߩu�VX�tF��;Xظj��I�C�3M��.��Â��j##�!b�:I��ֶ�}	`��db�!bl��;�(w5%�۵D��w' (V���2�R(0��ⵯS-̚"�T�V�e(��/��OZ��CXCs��1�e�õ9ݬP����Sn}��-��}���l�Vw��4�n.���Na�C�=@,O}{�Ȩ�k��^{2��o�Ԡ��)rX��W��O��Qd����-*ь��J���b�e��%����,G�Q�����?��K7�流}Pߓ��8�I��@Љ�����}�Ӭ��_e��[W	�����8�p�v�7Q�oc=���h����,+��RT��+ӕ�5r��P�`"?�,<;(O�@3u;�GGY��cX���ֈ�zՈ"��!
��N�:��28��i�^��͢$������Z7nW!(�N���<~Ќ�+F�J�nܟڦ���`��X�s^Q��_��!p�y0����"q�e�`n����g��~����z5H��ct��p��(x-����9�+�s�� ����n�?��Pê9�_͎����ݱl��e��l�3�ac���MoKP�c��ߊ�ݾz�W�&B'B���;Y�
{K����<����N_��Pz�k,���x���l^��i��zI n��3�z��G���m:�.r橋�UV�b5HG��.�I�Z��W)��Rx��< �/�׎2��IK��ʊ��#�������j1.;�D�}��75�/l:�;�gC��o D	Ǉqu}�(���l���J8+����c��O��[j0���ѣ���i	������k�_e�\����7�	�]P�|�W9��5�������;`�c+�qَ*�*�?����O�\ц�n;��}]�ZX_H�f���=�)z/�๸v����Y��E!lG�R�}�0c��5��G�;ND�O�qO��p&��+&��X�s��d�u�{�7i �V%'��A�H5��j�k�I�a���	}Ӯ�A���X���Q�8]_����Մ�:7�&a�,�	S������S_��h�`���8��*Z��S�r-N��G#�����s&��ƥ|��»��@s��P娣a��q������d��ٱ@͌��(u�0����LGc�b�u��QG=?#�I�
y���ku㢞��SJ]9M�CɷTޯ�Ύ����G�,�'�5p,[c�������+�mn��pt!�/�d�s�TB���'�NzF��u�/g:޳�6U�F��������=ـ�żսz�v@�P�K.�1(���-hu�vy%~��a���C�١��}��~G�P��$��A���jG��\I�-eە����@X|Q�3܇l'}�g�9��Z �T����S�]�_�0J�l0�e�hQn��X��E�~��l]�:y

�uC�TMp���y�}��'e	>]�9�� cz�=I�:k4�7A)������o���j���CZs>c0�&�W��-���(2������ǭ����5A�4����;��ڂ��&HOJT ���� Vc.l;�\���G<,�ihO����C;��N�t쪑� ��ٿ��ٜP� E�)�f�(�("&,F^�K��2)��@�i�,� ��n7j�[�O���#����@�?�{Jwy�%�p=X�9�=ٜe�D��ӆ��J٤�є�翚 �tqYk��wCx�IN*�Y$xe�4br��\Ъ��$�2�#�n��%�|�g���BEn����2h>*���&ܸ�ʠ��Zw˵�~+�q-�D�
X�\�8m�j!�������B(=�F�"1m�I8�2k>�7+n+4GDuejq�d�ʥ2��
�6�e!�tZpS6ѵ�J�!@�yn�W7&�N�7v}/�L}��N�c����0���hgUhYԾ�7�r�/���X����z ^\���>���nL���!���ǩ�f��Z�K63���PHF2�-�RW���o�TH�,��(ix�.� ���Z�Ꝋ�S���m�q��s�l�"x�~�����?�s��<�d凪$��FZ��k�r;K�GuM��pLx����H�[F���p�j�v��\\jP���ʎ�D6���cO�C���N�☪o�,%���x���5��t�����T�!yg��\��g�N#�@o,1.<���;�NϷ0�bq���*~D��	H3�4��!��:?Q��Sb�����R
���b4��%�Ɔexq<)l}��>�$���7k�gb���5W���'@jC�!2Y���	�
���O�`�K���Pvd���/kq�lp��8��AK6��N?�Z=��3��p0O:�;wE��!��9�F���M�g6��. �X�^�t��z^�G�������ZԙD�����{ʼr���&r߆�0�E	}�(C��ۂ�F~�Y��n�gL9���
����=��T��P?MK��[�$>�BǎT�c9F����>��T��"�����J?>y��Őt$u<Ʊ��d%ꍟ��r���D����cͲ֎0"��	�"6ec"��.G���%Y&��-f�ۗ��`љ^\P���hmt�����ے�<��b���wi~��o�Q��a[ɒx���3XA�λ ւ�D�ʈr��6c��̞kuPJ �r7 �A�;52�Wep/�H��r������l��Ř-K�O��`m�t9)J�:�ƾ��{���[_�����~τg��h�»	�B�� ����!���h���,���V}Ғ�rR ˪�YM�e�{��RKt�[���̊����EJG�hm���
n1tM����9٣�gQ�f��̲�T�����2�5C-�;rN���B�X�DeE�U%h8��8�Jهڟ���gM����P�퇟��x�N1�����4>�â��	R�=��Mi󢜑*��͜8�t�Kx� ��堦I�S|-�(2A9��M� ��9g/?���N��i���|Asf��!�,�yb���5z%o ��|�+U^�K�}�)�DxaIm��� �bIG�@���=ᓳ
yS�Un8(UD�(%��ou�J�+f@5Բ1e�8�$�(�N;�
g,V�Dl���+B�n&E�#.�'±�^�������59#z
�ME#�yf�&� �ӆ����O�kWF�xa�&	��ڻ��K�Q�����^��pœc��0�����\����pW$����ںE�V�h�5]���1�hwHu�m*}����{K�B�t8DE�3�f���t��NF!�������1��[�sgo]~�N�^fH�Gݙ�fՉ��<�O�DK��[����.�qa{�{��Ҿ�d�2�=�h�4��>�ۻn����#�9�$X�R/���.
�.��PO~�*&����c��-��Ÿ�i:3{��F���6J�F벸Z�}Lb��C� �4h��{���o���NT��E\�#h�_
"~)���C�*�i�voEޕ�<�d6A� 5�z���{��f»Z|L��Œ��\� �=İ���g�\����/���Vo��C~�f҇��0O,�98����$�m������HP��� �x��fW_��(��R'e9	�$����E��+���!�BY�)�y��)��`,,}���C������| �6�߳bKt"v�	) Q���#!�����f�T���bl�2D����j�R�"K��c�`��|ք=2O�$��񵂛�:]�DuE!l�/���VC�+C��~����2�,�qX��ח����۔���&a��J�f"�1�W?�)\j�|{ԩ��9��є�\�kH(�TƂe&�������[AA��bR�M� eW����/I�ޠ�:O)�%X��#&X�swf�Cf/��[��5�d�ʤ^�~��a�����9����k����"�����蓮D�?6��s�v^�� I����PJ�6��>Gy4#.�N�ɶ�������ǽ����M��?��M����߹��:�԰�\�����808�wgf��(����!���s�347��Ȗ��0R�Kߣ\$_&�o.	U��lR�c9��wc6�Rô���I������W	T�y�ߎ�k����Ŗbh!.c� R��N�	�Y���O�b\���S+A��W:ܘ�����o�q|�h$Q�Ȳ�k\�	K��9�B�nPc0@)��l�d��-�����{ f"J�u��RS��~�qɧ=V��9��b��;�/~����>"�|��7�ҡ���ӹfD��Eh�܏W��������bw\|9�4X|�)�-�S�x@$q�0���O|}�?X�%d���S�r��ƅ^��^�#�O'�A��e�;�����6�b�N��#>�$�$����G������W<���'���V�,�V�QЊV��MKv2D~�pŻ�9{�;�A�DS`w���Xd����
˧���7���¼QBxƙR��D���ٴ�-���xę�31��h�c}�yK�Bh � �-����b��?�Y��R�T4p)�Fa��Yܤ�h�m[�*O����ߔ�;:·�~������ *��S�`yJ�\�*wʉ~	@���-���S�blu]d1Q*8�@}E��I\�����P8֕�p!���0/�Lh�~ �؏���!�cD���p�I�'P��ks��G0q���@]��Y�����gb������$�k'������w@:��p��X�Bdw飠A����{yQ".�T9�0��Z���!�"ZӤ��^I�	�]Z��ǘK�YU��Z��M���}�%.�{��6��� � So��R6��2��L�����߄�!����;]�@yi�7O�"�ڑ�̸0e;�c����%挟�-�=��^� �����]���(\��yl��BU���� u���wd�N*"��0|?������ǚb�Z�t�.r���o������X�%�_������!����ਖ਼˻C�����S�AR���9�����>P|�s�#W����N�	����O��@s�:w��toI1��
��n�a�r�O�8j;zd[s�����Ӯ۷ݥ�"����J��H��U͜S�q��l��U��i<��1M��E���4u|��/�y%Q�n
>�̊��fP@�Z� 0��������3O�ONz9>[��V�_]s�4�����%n�T�:pP��P��מ�H"�����D7����~m�)3�g��M�G�o��z�Y��ɮ��@�({�`���r���T�&�,��`�*D�i�� �݈y��z��LN{��q!���-x���4��g+�N�b2�Th�h�F�y�S������6F�?�	l�1+��TS5��*��y����� �)�Lf�C2c��1���څ�9��v"+��̑�hsb-�����(��Ȋ�(�;<�����ǒy�EI�lg�2�f�q�P�ŶP��xl^�����tægI�0Ёh�<��+l	�j��Pl^��(͈G':�a�%x��Y�5�a���ڶ�/���:�����5�Y�I��E�˃���D2��	dv��*�_���3<��[�c�8��l[Èz����� Z�[Y�!�ȹ����kj~��K�� �5X�>�lZ���x���ʇ������7��*�[V���n��Ie��m�:�ڇ�8�+p��� ���-&�vuJ6J0۶�^���Qa�~�b��V�g�K=��vIm'��o�m2�@y�,�tb1I{��3u���Z��q�i^����M���~��&��$�A͋��N�="do��\$��H9����k�" �_�Z��T���@mO!T�	��2���u�*AS�9�w�rD����L�|��츅eb�TS��Qe��T��9�[O��}�m���ޓ��ئsѕ�=2�.B�1J��Dg!0&�K�cJu7Z`���U�>;1�*��c�-�T�6Xţ.-�mHpCq7ٰ�bQ(�7��t���l���V�9�c�裮��%�I�
n\1�����0��R:�K ��X@H�k�P����(8�xu	����dN�m��4$��M�`U��� p��hηӤ�:���Lj�=z^l}?П�2���"����.ڙ�k۾ih���.�n��jUu���f/ǆ[Y�>]�#Zy��OZ1r���o��Ƥ��^��P�C(r:Y��4���ܕ����� :X�N�3�&Dy�a�l�zL3���2�d��AL��Ǳ�T)Ac��b��M+��_(SV� D���d(���f�G_��6�����PtCsG�r�/qU��:�V��*�1��"��λ�T�'w�F*XKէ���;�mx';��I��>�ri�Ѓ�
@i�3D> �L�A_*��qD��|�j6R���UǍ�(�#Xc���-s�}�p�K��^�#jn.�~q+���ib�H�Ǭ�����"
_���Ēx��/��D��fl��,���Ky��#�&Rȋ�qy�4�����x�C,n'�W@L�}�M�6�?7ɟ`L��H{nl!.�������N�y�1�%�g��O���e�G~6�Kz9���1è����4q7߶g�*2p��@%�DaVƁ�*\,Q�G]ɯN���iq�	u�/K�Y��%�-	��+�
���@�7����!hY/�lL�y�\�!5L�w��������$�=�"�q�0-0@�5����P�fXv�>9�'=:�_�l-���&Vzz��~�[]���r8��/���t����
p̎�B��8h>��cFk��찌�G}~�ނl����^�[>��J�X�>!��\G[-p�s�}�:�2,�r���}-3�gw�|���'�za(9�5n����|27s��U�//Q�{\�rR��&��zOBѹ~�/�pް5���%��[���0wM���Ŕ��
m#�%Y?�p�G������bv���I���h"�bQ�Iɘh��]o�mׅ-��=6���$ӛ6����������uD��%�
B-�Ҟ��`K�x�uiC�W���`8ܫS�\6,�<���D*c#hކ\D���_�ZO�w-�2̦ !#��P��;���9�B���9*b�@��f�/2�[{�l�v_��9���`��L)
�c�9���-i) h�/Y�3�L66=}��]+"p�5k�*8��9�, v1m&��
�I��g����b��E�"5+Ы�kz� F��kž���"0����=d�����ʭw3Mfl^�+�v�����M���q��L�)�ݳ�OfM��r�MfVLA큅�V�D��5Ы�j�K���8Q���p�]q�_}@�`��&a�Q2��N����p��*����T�L�WP�g��Aj����W��c1s��ݾU�m'�I��f��ܔZ��a����c�=�S�7� _�º4@�>=�s��P�w��$�!D�O��R&��#��V��-�/�rHnr�1�?���"���5��Bq���;�B^�8��o1�ke���>����՛p@��&h�0�XW-�a')I�Ω-��6U�jK#�?�$�q\EzY��8 ���bs;�/�MKJx�/�u$�����Xg��z�d ��3�e}u��&oB���n�C��S�������>|�^�;��^��`ݡ��%�&G��~w�P�Fj�$�煺�Y�E�+D�0Ht{4)>��o�˴ƾX`�X���cT�悃�a����y��Վ�p�{6�3����y/�A�9�PD�^>���?���W/�TH�n�W�~_�$��8@X��ߚVi�$oۚ��n�� �����se�gK*�e��umat�r<�@س��؞������y��k��%��v��r�{Ȓ`"�D"/�8���~H�����A�AF���Dx�%�Z�Չ8��Ļ�>���Yv����<�aq���5��h.�����QY�L$np,bwQi�p7��d��/��R8�*�_�O���A��Ի�mV��L�*�ey�7��B���D6�3��`G���k>������ q��V��*6q�K��ʨ;zD���H5,�"��j����^�r�za��u��c:��pĜ'$���BS�w����ĭ�����+��:���D��)$ {#�uSqA��x�^���&?Ƈ1�p	B�\f
���Rg��Y`lУ^}L���Dc5l�]
t�l�gƾ�����m�R^��gjT��ee"r���Še�<uc�D����%�~�.����IIvU=~���W�4��B��\|��~R1,�P��#���b֔ITؼ���FH��6��i*��ħK ��į�	������[�nU I�+�F��`����<_�U�i���v���$ƃ���1��CE?q�"w��[s§���.�"cu3W_�<���z/��j��q���|�a"W�ͩ0!�8�/�#�[[�Z�}5��؟�Y��2��W�.4Fz^S�zF�����j�s�	�Q�BH�d6�۬���A���b��K6u5P
�R�pk;S*�A�zhO�[��r�Uo�P���X+c*sQ;d�8zk�(�6 ��-�R��b��N��3t�^��u�&�0��e.c����ԧVo�/� �{��A͞�r��lJ�/�G��w�_��y�d���5>�X�?LV�}r���G�r?}*��O-c��ja��?����<�Eex�'PE���ɩ���iy�Q�����4�Yg�.�W�LY�M��P�5o:�<��(3a��aX
��}��"W�9;�)��vݜ�/�>�NMj#���h���k!�����˔���c��D�}\!�s詗<��撻�.�[�,.���j�q\�Խ���]7�U��]T�� o���P�?����M}���
��o� �@�q�tH�l���90';��ӂ3�A��=Ƚ�/�d���	T������Q\R�P�L1�-��﨔��d0��z����-Յ�	ot��B#�H��)�u+,�� �0�\�z�/47���ߌYx/� 'TXt���^����S>,?x+�&�YP.�	��΅a�ee�I��8��r�+�/�~�Ln_�/��>��Oxk�wl��Х��qÝ�*�((;#�@æ�\�X��
���Ⱦ	��_�,K�d?B�R��Q��pO���ޓ��H�%M*.��CiЅ�)�3����dƪ ����Ef���;PR��W݁SqGs�U���z���2���ʁ89A��B�����'�e��N�K	���*T�m�M��RA��Q��%�F	��f�g�d6�lsзϖkpi�W��-frp��G��q��H�t=�LE��Q���e�#�!���_/�8Ť�K��g��_A��)� s�A��0I�g8o�+��
�%��>�A֔�N�ϋ@��"J^@�F�p�:߂Q{��§E�<�QQ���g��ᛪ�] ��o���\�V��J�R�6�/Eg�>u�
��3��t��,o/*�(�	V*)2����g '�AK�r�х"�sQ
����bx�ҡy	�����\곬� 2Ȭ�l�f�]�1~�JfLMD�7�����{�晬Js��z��L��s����@�PD �`I:��<�>�t=��9֙H���#���yx�U�O���^ ��?�G)5��Ҭ`ȱ䲐��|�Q���7�b$d����&C�W����\C�r������� �� i�A�gjt���#L/aS,$}��� ��H
Oҏ�|<��ecW�-xem2@7H��Y���N�t���{��9��+�D���ח8�z�.1hjIt�}��-���S��׸	`8V�fP�)Ԝ1��3�?�40���{�����p@�K���K�,;c�\rD��6t��w���Xfd������;����w.?�@@�D�+�8�v�(8m�T9`��(U&��y-j�΄�N��ΜG#�'��p�����=���ưr�?А���`�����>�~Z�=�,RT]��3gk���i�uN�sO���;�񦞠����;	��寔L-�%�n�S�Z�+A�E�`VqR0a��eD��-��z�ζ,�V;�6U �&/�ֈ(��#�Z��/���g���	�;>�(�t�ȴ
B���/���ɿ�	�@�b�����c!�8Z�08qƚi�P!�I��E�8�~�T�Ctu���C.F$	"f�iR������Ȉ�W��{rg%��Sg�R�4A`��|U7�*����#��<(�a���Ts�����PU�^���	)IOP﫶I8�������4�N�[�om.K�wy��(_����X�Ӌ��q��������� )��6(�l����,q�
23�5���Q�53�R%{�)�9��@M��#F��Sc|���Ѣ���@i�5ڂ���a�+�HA����"�7ˮαPu���c�{�J@My�iQ��\�[�!��y@cOl\>`|�C�'�̻�!�̉�`np��g)�E۟�Dy�Ǎ���_;E�_����ã�jwKݗ�:��C��n7�_Lz�тb{�L�D"��8i���	���(:oj�O�n%,?c;8�~��f5^���<T�D^���.G���t�V�1�1p���8��R���-�M%���A��"͖�Y����ӂ��A�g��UN�*\�\jٍ`@o�)�ϑcys(|���rT5ڐ��W�Lm;�Ci(��� ��P��P�zC��.;:������L��,��HurN<~��B� bg�ר	��hw.-_6x �9I��KJ�_�)����o��iN|��)y뷎n��O�"y<[L���^���2�ogN穂sCؗb�\�,"J����{09]���S��郔�y=�gwe�ɏ�� ���}���ʚ%��l�e��
���� ^v�%H�K]^�\b9~�x.����=���-��񂖯6%�O�Ph�SeQJ�3����Ў9UX=��s&
�L�.���A~�J$�U�& ����0�4��B��05�q!�#9cLL_ғY�A�t�mY�]��<C�R��.��E�{�S#�s,?t�ʳM��t��w���?�G���(��^�\}bV�$.�|Vjh��2R�YDX	j��4B3̦N�h�Q#�D�މ��F���E|]�RmO��(��L�@�R;�j( �Y�u�SC��4��Lfd�)��WJo����bT+/Pu�tȷ��C�w�*��~�`�>1R��	"(��y!�m�n�A@u�Q�.���^��f|v�K�������^�d��-��Ȟ�%�����m�p �C ������J�7�o�/ �<��Œ��^�µ��⺸Z[��o{�wm�;l���l��@�ىF߬��8">�27( �=V�1"'
*.E���8�`�
�7�K���w��J�%�&z;�����j��5�B�,�@����ʑ�+�+��M#1k2����%�)��t��E5^���7bl�N9W?aaf[ )���?�;K4Gn����"�=�BVҼ���� �U��8���}4n�)(kR�oc�5��F�|w�~��:��m��<|>������W:W��T��(��Mpd�"y	D�/^�H+�8�A �I*=���t����FC	�n���m��|������[�vT���K�Ps�N)6\� :ts͞`�����s��r[��'�>���M�>;�Hp���%a�q
�J�y.	'����H������8J��-(	�4�8	����T@�4�T�dy)8��t���]���+c����q�i%��gDL8�$!�3���q�g��K������zV�'.���M�]�a٢eh ���ia���<Ė�I�Kaw��G�u�Vz�����<7���4*)��Փ��������p��w��;H�Ũ�bæ�@�m�"aİy��g>_o�S���Wj�k?v�{�{C;�@[��zX�"� @S�4 |JO�1���!8����,�mʎ̹N���nT�d�Lw�J1��l��b���\�|~>�}|��Zc,�08R�+Đ4�Ϡ4��c��ʈ��Y��ŏ��!#��\�x�q�j��*��%	Dn,GU1�3n�~�PG(.�MI@/ZԌ+��
�������I��}�޸�uW�b��cU��8t��
%s蠚*^��d	SA��L@�%�� �����R=�céVև�D�%ċ�l��yw�Цs�xB�M��Xǲ�8����|NGF�J}pW��%y�'�]�u��L_�U�e 	!��¿�٨�)F&�ڇ柢Ͼމ	+�1n3���AGo��Y��[t�ݖ|�wmz?��`��X��?=7dzf�@���푍!��3�Q�Ȧj�m��!��%��~[8���3O�k%�5�*;U�'�q�1 �\׉���� ��P���(�U�z=`ƥg�gֲ�p�gj�SsF%�)� y% x�j2�e�|b-r��?��Q2&;>��Ƭ��t{�a�bZyxn?|C"��h$����rJt���i���]
� $0��)~�o}���7V���*��j��dP{:��\�J��<2g�oUh�?3�F�F�2��'pg�[0>F6�҆�6��+6S��ڴ�u)WT�y�
�VB&�^�B��J`ky����b��c	M��W����J�-����0�f�_�������o mZ- �P_y����#��<L���i�?Dt@�i1r��%�u� [-:6���W���uA�T��U����b3˰����3�g�F�q�6=%]I%�	����\!��q�� �������/\��#��-Ȩp�X ؚT"�`g{�'�)4�N����P��q�� ?��C|�� o�L���6����J� ^�ޭL�ǡ�84�|��.�!ϖe�0)�q`[D{�'ݳ���+�6�.>������S���J1g��8��Q| ��&��A1 �����'�:�i.���&B�`�~�2j�9a�����K�9��b91p.(������N� 3�
���3���j��}�G㲥b뮙���+<�zet=`hq�Cq����o�e������-�1���u�}BR������0"�}�� ��|C� �H�ҷ�g�؅�6-��ˆҫ&�tʉ�Q�m�[�?l>��@�rE]5`�Y�� �c��D�׿H^I�Hv����܉%K����Ql��&�°��J�]�7��z�~���7��yYB���DKgc���^�M~������)DM5��?e���l^a,����wi��@C2�-#����@�O�0ρ�?�F�V-�Q�?���%�@{gF��0���a�r^O�4�-��.�Ƀ����IAnn���@��_��}��� az��
�S���)�M5��͙�ü,��Ҡ��M h��nو��B�qt�|����A���Z���^W2?/�u4���
n�g��~�B��)C���D��	4/R~�̹
IB,�y�Cqm� ��7$TwJ�U�+��!������i�;x��EVX�E?�IcI�;k+k���|d�x.�(��a��<�|_\~1,�c�����O.�tig�~v	��י��\z�d�V#7܋d=�w��nb�>K�\*d薪��ա*!�c�H��$-'f��o�+_'�6p]����v�|����ew|���f��V_�Sl��"����)>�sk�Z�^J��ɧ���ʏ���n��E��#���4���rx�V�ĸ�4k�RN^���Yc��'��_�N��+�K&����ܰO-��O�i�/SAAL�ki�t4�m���
"2����.#�vk<�T���Ј��g~����"�l3rj���+�8�D�d���<4�h/a�2��*��Π����۪�j��l�u��ˊ����b� cًz��S@��d�X	}������P���oP�d�͑��y�\lIrJ�2;Y��f���K�<E�3!s��̔o��O�.��f�vPt�0\�z8��<��F��H�<����^X�{#��4�J��5f�M�D��,�dGk�ԇ4
�0���揥|��9:�:�XvFH<F�<  1 �]&�ȖN���B9&E���پ:!�iR�"���4�@s���`���\&$3*\�&�MsN���y�S��J�hV/^�^3W��3��_���ҽ��B�������	Ҹ���e�B@LdZ�y����Ɉ�^��=M3:4�s5F��v�
S)��ѭ��~꼸�1H�	�~f��r:2�/�Z�K��j�x-*[mU`e��C�o���(B�6ZV�>�e��� j��ל#I]F[��şhy\O�>X��S �?
��3�d��w�ת��ă�g��.���%��+ʢX�si�L-a��WP�j���9u ��� K ��j�̼��Nګ�������N�eT��PzC=�.+&}Y\/J;Z-�I?�3⧜X�<D�x�zQ	mNR���
��� ֨��Z�,ӑ����W��4�=�-k�*�����I�fH��f� �5��.�OǑ��2�qʚ���ct��@�t"<c������t-V���x����$��^��l+�Q22��pk��(Fh�R���b���i�������'1m0t�Cm,l`� �'yB��O�B���̑1c��R�����zvV�[/6./�����p�^\�ϰ���+Og���ٸ&*�J�-����9�;aOK�����E����=Pe1%uG'�H�<G�v��po�L/S����]Z�Ј�C�]+�K�z�`�O��\�D���X���b8����[�b�(4̮��d����P�
A���DT#�0��;E����4�ƥ|�sk3��X��1פ@�Y������B	�1��V�|p���N�m�yET�*Is�n�e=O{���J�t�	��tJ�{U�a��?���6&O�ns��E}É���>����u�ō~Ʈ�^H�s��Eˬ�����Pˀ�܌:JF�{�2��ID	�&�`&x��O���K"�BP�xmS�?>�
PV�1����j;ĄE� �W|C3S-�2���MWn� ����684y!MK`(rz)��$Gk�!�X+'�e��N�~�6� �����
蓙��[<e��&��<x=��i�r �e����{D��Y*w�0�8c���^f��E�%0�
���ZE"��� S	l�g)�.��C9ay��=d�2���0�����.�������>�]�r��&a2#�r#|~��~�g��eOڹ��qw�=-��a�f��z��Y��#�������A�eUN�cZ\�4�}�п�����Y��m���Ňy���Q�GV��� ��2��8�6(�����9@�����J-E����$�مR�x�3l�>��}�mN�Qy���0L�)z���OR��H����r�4ތɺ���?��7�=���%�,��;�6X���+��7��+���.��'E4� ժN~ʛe�I�^0�NRU�5����{9�	Ѿ�ܼ&�akǷ����}�if~WrH��k�����7A���6�f����cQ�ɘY�zӕxL)IyӒ� Gb� �D%�{����CYdu���#8<��uE���Ѧ-r��� �	¥0�ֆ7��R2D�݈���z^�
$�T/��Y\�%;˪��}f뙐��7��i����FqZ��4�kC�^���Jb8iT嬼�N=���GD�p�v�Iw��p��6�<�?�������� �%[�j��`����)(���E�����4`��9_@�Bl�J	ɵX!Um��ˤ5�:ϳ�:��F� ^���n0�no�?.�mg<2v�7��W��#&[�s%i��r�j��2�l'f�Lɡa�POX��)��Q<���>��>r�?�X��-r��Mz�iF��[f��Wb/҅�[�	܄Rr4�.{t�Os��m������kM��.h��J��
 F%▭����h%$u�pq����K���]���J��_M���}SZ�0���C(��H%j�2�.�¡��~Lj>)��u=hi��<�����Q׎*�z���,^?ܷ��'��Q�j<8��9�wb_q�9����]W�8*S\���u��C�+����z��ӫ����[�T��'F���+�q�#Y?�Qa?�k����<�m^�[�+�Q<�CK�&<�#N{/��:��F��
D{���ro/�lhE�+���B������U��H(:{o��_��u�8\�p�[��\������xN=������zy'�qY�����yF�}�ҡ�z���w�ea��-��]��ku�%K�-|�&�b�G�ĳ���I�Ӡ'E:G��Ly�����`�o��f �E����N�ҡY+&��V�
jq�^#�>��$��}� c�W��5��%���T�ڀڄ�JM}]M�P�Z�y
Ye�Pf�#�d��bu�szk9)?�g��vF�qA��[�@Xv�alZ{� �^w��b�s4cs�c�~��z�@�����y7d�������1�HzL�� �M{������38(���H����Pt�yC�:]��\Oh���/��wT���Pv�eX��[r���4*+�8�6ER�҄Obkg�9�u|����/��X^���0�v���&�]�79��p�1��4�ߧ�W{�95�;Б�۝��E}�(�b"Pw�d�o���.��N�f���Y��yVK�ѕ��HA����,c��\ָ|�{�:��!�͒p�h��R~�ڙ���JU���#�Jc&Ԋ�w�'��]{Z��8�9-��QZL�U�~%}�f�y�,d�t�H���\=����D�턛f8wF�X_�L���x�4��eW���r�d���@�D�"�#�L2�vm6k|�{�)=j�ZWa��qsR�M7]��j]\u��Z���)��
be܎TCҮ�%E��i���VCk��2�S�.�Ƣ(�eV=��K�y���l�}�D�#l�p����ξ�\��HI�0�Zt�s�;��'Ï2*)p�~�p4�m'8�/W���� ��c3�u!`��A�X.�I��hq�T�zJ��D�ܹ�̕@pEej�۴p&SV�zL�ߛ�=��5��?ʅ40F��ks�l(�x>�-����Rn�_�$g'-��'���F�Y�I؛��PT�
���;��N�m�u�SL�����oq��C?�l�Eb��;�iq�8��r^f+��{�S�*M�6?�:�4<K`���E��.̀�uT��^�G}��6�60۰!��zLU�� jD�8b���~���vѽT��@�O��C� 7���09X����o��E����g]�Ͽ���	{�2�7erj��Q�7@�,��g)�ձԩ	�v$�-����"����K����/��w��*y�[�X�˦@r��#��rC��܄&u��;���`���z��\���H��d��A}�["'�鞨R~��_n�!ڰ�H�m֒��B���`��+��cĭ�Q	7(M��x}��k�Q�_[��B�C��U�S7�HUݨ�d������>��fQF�$�O�[���ܝP�`rO��<y���<u�����"�%�!�,򭜏�h_Xvx̧�O�� q$*\c��<6����]x $=����Q2Be��.����ٝR5}H-������Y�N���
ԃ $�Sd�����а0�k�c�]_����^vOҙ�p��M�Ǖ�Q��Z>=w�����X���:?*���خ���9]�|Z�m�ю?Ϭl*,����3�)Z|�gIa ��y��9�Sp�0�hKʪ��b<��m���A%��Y����p^���6�ن��ӝ��m)�(��
_�~�'��iSm��g������yr�p°�z�Y�Ϛঊ�>�疻:�aL:��8&CcK��_�w���,�!����*=�@6��?\�\��ܮ���K;��Ny�%[!rt�g�����+�@���7_��,]��L$�+ZTڑ��Ŷ?��/vg�e���U�Vs��d �`+̲���3Ϗ.I���3;�s�A���ģZ֏!E��G�.W�c���-�8��96�S��T?����eJĔj��~l�h�hB��ɖ|7���f]ʞ *7�qm�z�C/?������漏�Udd]�3^�i�RI�	+:���G�x���C�H�в�+~�U��q\��,��fH!F��,�(�:�Kd�n��t��AyƱ�q30�q�A���|�v��q���^<)�����刲�k(�s&ꡐ4������D�[u��G�q��#<�٬ w���򉷰��M/F�Mѷ��p-Oi����T:Og&�B��5��d솳�tϠ�kKDX�`$K���c��tu�0����Ĺd�j霉��(��&m9��3Z��1�79xC�:��а�x7{N�X����{v�e1B߆�O�meZ4���w
���'�~0� ߎt0�6�qA!V�J�
Xĩ�'��pp�V�.�%�����{4�!�*�������Q���G���qNǃ�hwQJŞS���L�ܣԐ���n_P�,����I���K��
}	��ƘbI0��K�Z~���am2�V����Sܵ`AX9
m���1	���T"9I�]V��������\Cc;_z���d��K�]l":o��AW�a�C��p��frZ���z�."��#�B�׊0�e�]����*o�e��SIp1��h yӜl9�Ha�,�}���FRϝ�`7��ɋ1�GrJ�˕��E|�K��b��A�s;���,c|(CMa�kj}ϼ���!�6A��f��`%s�b��2/���fG++j\��C*&���砲���>�?�nE��!��(w){���{^���1�УAD[
�3��=D�f.<��8P�@Ԗ�*�q��"��08 �9h�̘p;�l�Չ�b��!ɖ1���>مQ��E1N�E۵m�$Y���;��B��!Z%%}�U�K(#C��t?�l�7��{5�R����6�!��߁�Y���]��;DD��Zz����ޫ6ρ�bЄ�)F�w�gG_W2.�����X_��W�(0���sA����Gb�1���>�^��A���F*�e�	�Rm�3�y���5�<�S��[�0�7��q#��~7�I�M�����E�������=!�Ĉ 1!�t����d4�H�(�_FVd�/���eG�`)�P��@�[�~&���b��� �#q����_���#b���(�h{|3R&A_��]�ʈ����8%M���>�L���yv+d.�s��%7��&~��h�����q�]����_��JŦ�UP�AL�w]�6