// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
iBNcU7yAWPGY/8GP1KAr8FxasnBM0jR1izEAnwBIxVdarFTw60IqU+M0rp8dh3Vict+iRGKlHHQw
WPMoy+X1jNEVHdWVb6Ic7g9732Enhsb3dOHeV5TLPTSIkJbjHOk38Sz43DcyPfhkdp/Nex0Xga5R
QlY/wNyOdtKZbtzBRB5DsDNODQhGW/BXr2ZLRvcfpq0x6UgcYf0VUqZf6UWoNOyGEVSHcNG9UvPk
k8OxWsmEqKGxgNdOZ4uDOuRg/4UBIBy4MOe4Q283HUaHu72lLEANU73pIBEy0pMbNcDGw5G8GJwt
o2J2jMl+01KzU51yMc68FsJ85sFbDzNnjNdVGQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 39472)
CNeFmQB63aQIzWv995pXCR3aL/YMinI0SGzTu3z+7ZOOU0z8DELtchF2iiFK8t6eGKrTTfBR/CUv
aR2UlmNnwo1pi8ueOLT42Bz3VIjGHZ48CppmsFisWhGfx1RXa5KgCcPWyqWIRo7M7SDJMuEJMu39
4iKF0JpPqtCAbWoz/zMVZ/2cY2uXynJ22PjNJ9G6plg1RzOCSSJKqopIknZUOmDsWv9H4UBXXROI
AM4S/P0ZnPu64A2DVTUvS6jvXGLxHxTmekB0m8P1hqvxOi/q8quB+QIYiwfgQLFI/bYXHDq/aetU
PqyL/FBG2NsvXJHYm/BZYtOj4MRd331qCpr1AIgRt6VvRBorQZEBAhiuiwkzXluRWBQ3aBw9p4Bc
8y2ebVGVcEfoh3fVnMYuOk/R70/qRRiXz6zvKMSKWMyyb3R5cu0ELxT37xr9cyRCUhs3sroRYM5v
UE5pq2Bsl8Ys/oFo7+NcZaCvQjicqPzDEc/f3uEymUBbCvLL637ylZmPEhngE7mlQzTGdTIjkyzE
8pRRv+xLobteKjG9iKnNRllkV9lZk8Ux7OIaFlv+b3IlaVHwh/28ZQiCy1zJET6GOX+Y+WZVKCrM
e1eVBvv1YzMyuI75SDOfuUcwX2VbzhcWmfi4gQV8DkHnniGU0H+UVSklhvmXWAvE3v+ActAgPOK8
B2qr8/7W/9LvGmBnP+bgv3JA4wVGHLxHrCZqryHTqcZpF6FAfr78uFALUnf0wIpokdIZAKztGT38
PttQWBds+VcDPsWmx29+sRkABD0ldaxLICiQ0yBXOagsmwIBqmzyhcP9XVbbWcyd/jojM6X+O/dT
/WmeVz0PbyNF5mDanK2c4HlRI6BR0ZQ0NSJXdVYV1U9J8XqsiXUC6/QHAqMlqXXui4TpSG4B5DPf
0Yfy4lFM0WtoEjPLHB7LmbQvouzfo/UpPw8oZFUmPp1VlWr7/k2bABWDhcvww8SzB7cOE4+bPnFr
eYUmKjwdn2wHcPgLJ9gWSRGKiXVilvkS4MjgTA4BO/ahc0EPAfCL/F3wdrfQCKvw97gIESAjwVyH
LSAeyvjq7p/83kT6n3pkqm22MXOKY7rz1qp1/he98HobqSI+SBhm9r+8PcTBMVSjvOA9qXTy10Qn
TxwjeSBUI144QPapjMdVbXUK5gKnl8H6blH5rJFNVtVZ40dDxMzOSLeoHK/AdCBPQij2NQqEGidV
5ymSGFKUGoh/PbokMA5MLueFJF1GPko7kxDItDQMFlJ01LZ1OROIBBTyqQm1fzzjl8tQuubwC1Kr
hDnKP7bakh1Ht1p/ariRVYCu3Yugwum+6FTIVcVytVq5osaOKD5Vw9nrgPiJQJ9hP5wMrfYThG3n
A/GJupJPHVP1QqqChOL7okaPX2M16AU8ccAFy3+9AUWLc+CJVs5i6yuWu9P+N0Dzsu5/Hce1iktd
lDD67f4wa0OVv76YRdBCT/zpaRYRnjoSyhM9dj1L3nbLPCfOyr9ar2DXrhiC2q01ik1Dqu+oyiNB
wHc1MUyaMuyE2D9Nc1QAFLUZPsWndERObfbR2SMxTqBS6BEuiCTx2mvw4kWTrUs/q0e9OKLe1Xvz
X9R5JLejxnJ3M7hUh1O/Iz6YAwSpmCzAXfH/EK2sNhSx8/zc5T4fmqnY9iVnbslVu9H0l2M+KBe0
9cQB+nztgtEr4OHGMrt3kT+xq+gi/PK027YDjclV4Jo5lrl5cLKJfWddLa9uGrDMgrNZZwnKVITO
3JI3dhoNu3lbihKN9v+jpLm5DN8bfRFQzHwP9U191U/+g/Ok6UBn4jAUx2QWh59m5F5I5yqYW2k2
cS1I9IwRamteuwPja83exb9u6uast+xR5KurvG9SRWCOuYddZQoKeMDDRLKwabRP6jw8a39a+fhQ
EyJYLDlIVE9sJitYjruNmB2S4XL8GW4vu0u8bjoZC7Darssb/9RqAZoMpW2IYWH7kxLAPTL1XhOi
kWx00UOSpIdHcgrRBwucBuUa9Iyoe5CjitkECLgh2uFO2OIQ0aRuA/Ej7nGTgI+fGmGefAn+GMBG
DcErc1L8M6dn2epWPqJwjjL4br61dTwPnceyAWZe7llMsZXCMEiWlwC/J0NzxLbTlsTgOqhWpd3e
IzWIz1pgENxv89rw8B0z2WHj/U8amif0mZN0E+Ko36ul/nXi5fLOiwktxiyYsCfDFphUnJl8F1fe
bX27SL7RD6kPGyzIrnsIf6AafxLu89PgwF0A9HqqmEMLTwobP9Rlv4u+bTPgFjQ4L7Pes4fB0ZAR
rOiuvoclrvRMbLOJQ0WlqZPN7MUeExCRfHE9IWeBZPXNSVP2oXatb3Ro1duINyAK4duhaNU1lVej
UdrsTBTUBVh772HtES04reLwr4oYqW6fESY5ngsZslFr5RVtmTwdmx62pPu6pjdV2QZl07qXSv4W
DpEG0ijqmu/u4zpJf3Ssk4qilvbyNdde4ivE1odWxLvdA+waT1tHcS6BNTUELPt0h+wz//pBK5HU
Sri662k2rsk3hvI7CsL12bjVQkpyprwJZ/2y/u3m1Lm2qNeiC+1MNoNto4+3eiQTJ+pKTf7k1hEd
NjHsmBPZftmyesXGeQY6qyuIqZMURBWPBSrHwk1mnGJtOBQ9xq9GeEhgr+UvZH05sX3fqMDeJajM
WDl+nK8vrm2ZcSoZInQnmjy/bhM4RGqqNEwusbDuZkytkavhCD9MaU+ak++kIu1o46H2Ecx5xxqs
0844TEyPX0pXpN8SA3VYlMq0W7qrS3VL1ZT4Wve5EUG5s22xWb4QZjg/exo1m23v3LLNoiT5VqxN
/0OvUNPbIcO32zYjJLA2OuYUNocPzGoX8KQFW4CfSUgrl7wg3qQzGyoocAkS42UZac0MB+Y1iN7S
NuyREVTBJbUSBRN3vhIFI5HGkbGC3IGOvA695J5xzA8LJpzfsVrUG5tiZiw2+5qnXQhLpUrVz4uD
DJrX+CxlVA7nWXLMkIjTtfH7gdwSnEQqRdjQ+tDjvFvI9WrsvAf+8MlDtlmbs1y9Ms/hlR69xQ7B
By0IIy3b5dBHI5WmrTwkKW/FdMFAd0Bi32/LNk4Fl8sdX2y3nTjeFS8jVodn6mfzOLPOaPjaJ8HT
Xz8XOJL6lKdXPNj9Wy0xX13jyP2XssGVeqi/B3yx7B48pMkLvkEGFpJ0+3IEFW9Ezdn1IN6DnGBa
VA8wfH50Bicq4Abubrz//VlbxOuoXkclnPlhtm8UrlLTFdbtOu8UGUWbQKSKcZfMWIBsj44IGE+c
llbrD+9H+SLfrCpNCtDIvBSZjwcF+HOBiciDNYyDCxzQKsMrKlXYp3RMnYYGNrzc/hwaDsYgPlfg
mGF3VeqLHYYotqCryACtIaeNi8UD4ZBk8Q9pO8Cpr6d+t0yQxDcUeh2hzMxqE2lCQnKMlmDArG9p
XaPIem5AAwySQKa0B64t3cSF/3ESUR7g9co7JEd6Qp/DpPzxQ8y+ytDzpUnuVeVqgsgNurveJKe/
+Eq+ygN0LKu+qS98W3Mn4Zu7/Yf5O1j+gJR1TWVBbF2LD+8KgUJhXfy87CJR2v1V44Vh20EZz5hR
nxFVvb+ElfYjuR517STFVcof1J86ZJY3OHAMIKa8J0sGI2DJ2iUNMfLaYLxQaJTVnqC3LdsEAOhW
aZON98Ft1oc7wE2ONkdvzgZksILM05hbUJxsynZ6i1NPWs8GHXPafDvarFydwxPJdyO6YMXBMZhC
GHbYFbXmvbPNm9Y5hB3McxqcdHpvXoLFJZb/CJ0BvPEEbMUbl26zUR8LHeIzMwAMZmg673S+0pPD
jJejY3sBV+rhoMqbslGAKOPsBsur4w4ytvcCzewE+4OWCX46BrCyqr4131yc8VE5YTiLnFTy7EFU
QAIBY7/YI23fAfktrPEK8V4ONsIv40gLn4ZZYUmTm2JYivmv7sjZblkU9D3uxMIeYKDLZu0ZrqXO
hyrCEmsqUYS9h0rbbJITyXdh7WsViAAZOzGKRNT4ShNeUGTGvwzoFcgUtI4tx4/667q4X/zPgn4U
QezWP8MgeRy2fkM92NgOxYAHOJ4nWA7VBe9h0uVuZipWWUJho/Btqk42ivHCl3KX9+2A7AZMpUcx
11fYB+Aqr3Ze81E+D35waSPtexY5Me4QYQQay9uDqU1yIQ6WK7FXREX6dv3OKI+j8nYFe9JUTE6k
rlJtdoteOih5RN4ji0d9UwMPedISZROOSTyaJXOJynHx2Wx6ZmQo5nmwvPP/PenBa84qNVB6A+aM
eS0xoTlvNmLalvCCE62snhYDKMVpj/BnjoAd0U3ia9++s1/KCqFmUloE5rwcAIRF/9VAop1XGKAO
oucHEFB3tHYOnpwBZlI9+bWYj91YSgBC0nQhygTZGXt5XrUy5AmXiWamDyjBQ47aXZ7nkZEE/Obw
/RIdQdCMRXwajMrxwj6dzYFDzYmc11JkIfmbVhbuVHWu17oN4l6reNUUjsTB4EuYEqCEETNHelcL
HdBaqgEK1kbh59ur+NEF89EkJptY7QcyKZf4YIdlHXvCj8+iRKprxA9JNynyLSRNc9yWk2kGGuvD
Ld5LWLkxpQh9X1dGmoACygOC7EF3kX8nxZ0bMelVw5BRrx6LVSiD+bFNCop1gd25onhM24YJQR22
olDRR6SxrMQBpG61+ztRsW/Sjy07V/rJ6uwxVt8R9zehsoljyfdvP80QFFTW8FUbfyq6X90XmFlj
x1rifKRCbr0vW+KjmNrMWiaSzycqfOC87GLCGlxqT4sDSrj+yk7bITwxuSa5QyRLAfhzui0FMZqZ
FmYe4si8YYaPjqh43EM/WvGmXqXKQUZtz2IrZ3WyRrnyYE5vEgAyeKxYRK80vgG1HNM8IsqKVtmu
5SnsQDb8cXD28mmAR1XpU1dultpoiVKDzZpi2OdGXIamkfSOnU/m8QZL47p01r/5ph8v0941cwdB
lgyVDP4y3FiiPHCXImmlcONAbcNHzy9ldRwF3gJsj7X/tEDsCf+g8h57xPe65bTgAC85oD8C1ULn
b6K4/OwDOL4MzLo47EmkbRnCBaLMaVffYOBrTleWzW0l5A15Ldfr3YLuMQIWViGjF5NGPDMGVEti
zka/kqUbuPDxlzMENzVWMN4KXeNdSwojViN7SLz5kq0UXlSxLCrNNlcMIF+Xd3Fd7yNy58Ruq89G
vfO4jxXQiuUs1KL9Us/yYi4AUAjvqa3Mwa1OZdaEapfkgoK9WGQW3pclC8Dytxs3VkLArJfuMnkR
o2JduPT9amguS9kwHZZRp1qh1zLj5PY1A+0ha/x4aZ/f0dQK4n5mWFupsseDZRTQuCNh8L4xQFRJ
W9Ggryj9+e8IAaBNjD9SkTNr2Zi5KJuBm3wSgeS6QQVwgVOu4nRlkrIji7ENj+Znv+b/sRzVSprM
gZYGjrtKl7oZe5QOQGrsewYlFNlCdec4jAVSD9eDsic14BSGKBt7hxDCOIqDN+GbTrZHTpjMH44h
ex6l1VoVv7nvHoAJP9nYYYaVRXBjtBykoeCVbdZ3Y7uEXZUzzxO6ZU7qgDjxJVr4DFIpKSbiP3ub
WZq3/J3Wxz5MrZ7eEG8Sm/8St/U+RuUiEaBW5aIKNwPHFFcHuiD6JMTlbJbRaffrBoQaao7TZpx9
t26djXcOWOMWRCo3HjvybOUaWFGWd99GYeeGHJh2HDujVLhKjx1eHvO9Zymk4Aicyl979jAkKab9
CvYGARPFtZfi98eSNMWUuYjsrRoAcQgsizc18Ew78QnsM1ivbxLOpfU1NObNDZXFwghpeYy6uQZm
P0LSiSZFVa88hr5lwXOmLgs8S+4S2MTtILdIVML6HawPLY6TmRP0+xed1YQi9cdAOYHHV+4FmO3D
gizXHeateDj5rXKQE+qtEkh4zxoe9S0vFKcHZt+d0UHiuSrjKUNVkgwL9BfIUypVccgei37QokRA
jm+vz32kxlGw1Owuko9XcVOFdYwuEzyUZN5QZebYixE69JbJao7EUljT4yz0ZO7mv91EMN0ufLPJ
NThBpbZkyDTvrwf7+fJhiktwmSr4nCdg8n4sQJLkRhiHxkYTCD/IBFmtievkjx9Jb325La3jw+HK
jMleNhD0sAbnaid2/CB+OPbv+mbsDk3dwM73I8cjcCA9ljKgD1XwODF11Kl8kJ+JeazL4tMeLJnP
cKsscKE6Cg3sbh0H7KW8IzEN1RTr253qnequPBYnirA8TxDL//qzDU3o303xqmz0gCNLUHxePwB7
diha7MKlbEYnP9xcbexFSQuCBLBqa3HGI2AbY4zkUMWnYoorENhym00P0B4yAsW1ivqdrV5WBeBU
GV/pqmh0n/wS6ld+/GQUMW4OR0yaaISI62p5FKKPcoUSUDqRbjoG5YzO5XjFAh/fPxW75Wp6XNz9
BRICJ/OyHZNhZQrBA2r+PR1BjDM6Zgal7b9kjOI/8JkuC1cJ4BCEL+/hmsyZmHar76BXm7LbAo2D
epQHXrhB+w79G2hZ0pj7iVs47gxmqL10YGcb6GEXs+lK18g94i8ayBJ9c8+Tr72Lb0A0QT9BA2B/
FtXfjZyZzAKeimrgJR1JhgMHqNNnKQ0eG+GqMCgpZknscZ6n5G29k5poROHYrDSazLmKq4j3KcgT
CpC7ghqIIXftAp9depRlOwWBWpBk8MsJPqnCt8RK/iBDy0oxm+aJ8gojd2CpmD5VfSZGtWdxP4QE
gS4vkqKuaWWlNt3gItMkbCfj9gC6p5VeWwz+J6FAjn3s281UoGutDVbKQzYM7B3ksv/rC7XvpreG
Wd+wmC9uihB/NrJbkr133kPH7DJsgT/29LK3bdb/Ypu5zXG6bc1QmrXjrDw0kfllaD3zMNgsEIs8
vWs5aJPpxQUjWQ3DWjAu0It/SfePDQy3UstTJ3TRQ04nVyzxdn8ESfcu9ktHxIwFsDh1SOln1v23
v/uyoH5FWAkecOobo5w/sp8bJeIP9qTSbrp7zooOg7mUcopHjv0VasV5Gnh5Qq4OcF1xhFpfFpuh
tLKTm2pDM/OdhAdqc7BPZUdJ0Bz/YV6ss2Dux2sgoJGHwa7Ocanpu2eTfDLoKbm56zlNMlIbrqSh
9LNXHWPnYt8PmXJomyp+D1hrueOwVpIMXUWUpZF4snpOvduxIGLtHVdTy6T0vR6niZbkE/R6CnwJ
MudCIo/mqN0NzKtaRiM1rm4SfdV7+PA4J5QTxWheoQ6E/EstvXIeM1/laVsPfHKkzrIAp4AROWl3
/TJfSA8dgzu2Fe0IdVv8VtAGjfIthAQOf0zu4DtbQvejxNjTRtw72thev7OX5cfyFQDQchW8LBXA
LX+aMfiDX78V3d/wVGAaawd9eh9RdmtHqjc9bp+g82o/UQEM+TYVxEsQfv77ucGOBTG8VZRiAc6y
w6xM5RdrpkwDqn7mz8LpNxw+szpF4gzWSkqxODwaLfaMQn/ViRuPXScq265QENpCavPq4pc+5xmk
fhpZmgaRyDhbhvkFIw15cNywVnxgnUEzAUlHRSm8ocKCqYiHVbDZUU+Lo5uDnRtWGj8VPil8TLvj
i8SQdXAyfrbaIgo0yTWKsntZDU/sOKym/viaaqy7wfsSj7r1epAMkFjA849odCOYG/BRvFHZ0Prr
5J/8zeOdRQcgoxEzjUxz5iuDzXaXkBTHxxMMWzwtoD2HVcsHIY132lycag7OVNK8IoU4ZoUiMZmV
SDfsl4HsjUKOtcAK3gQBlmw0Q1swqDmtDgoqETG8LenYhDNJZ8q9gEu1hDoX+0lPoipqO0CCx7UN
eJenElX9kmVJK5Fn/EhZYKiEjFFojlW60efX8ZGedoIrRIcVrpj7wEOl8CpesWFxQ/Smw6tfJmdx
XXhucJeUN3Ys+TNEZT7rzqdFGtdQJU8FVLPD51XVMTMt0a6Ej7d6i+rK4AdN4MdrEZQatdpWXVCI
05r1bocNYxJYfX2TGayr6T4MJCFB7C5uE67Zls/vjRRKpZE3gKwc0cHpSqgaA0r7ChK9rqEBpveS
cbD5txGABs9uB80PD08St9UsMxsQUqU9GemQISUpK0rB7UnNn7eusinw9DCsKIHspHLlAGpWzwP4
FU0yFKm35v4RSOu5Ai5kwEJMo2jmtcNcVHXmRK3iW0w589EhMMtKl8zw7aNSudd5Pb+24auWemrG
FQXN9i+ubPh+/WEZlPJgG2ppSnjyEtCBb8euH/dodwkh2IoJfSjgKUM5jltx1uZgL7WSmFyIXl/Q
Gy1sF9nnbJH8o0cmbxjbmtA+YZjJKAwTzKAv69sKZfSggh+y/Ik2LzAo06vFTnX+KG1oZs//Uk8a
6VDjMAhi+qzyYy1qbCRioqm/qgjVrMQldZUVpcfCq32Ugw8LLLK0UF+6IROOvcyI1G52Keb50cgx
KggbP+zlp6qvYo3cBIghFKTQ8SgD4MvLYtCjN5EjCpjCK6SftMQ7A0Vq+mKbMYHDImNucPKfIFkv
z2rWcqh0hJSQUV7MRCcTJLr1p6TKTYC+nOpFZkAeQ0VYP06hrSXhKpdnoyrSHblzw8oCVLkmg/Xb
pGfC8GQ4+Fbfait2yKBcKmplTS9OMeuNsp320OsEqOkg8FZtvl7Ox3RFeH7DrX3J/pY8ByIYxgy8
OhDamlrTqjAuflAJznnUTPqujR3vHzyDE0hPZuZ3t2pnp1ij1Z6cEJLFNmLN2GRshuVOPUFKFKjK
bqJ4G9yc/6Q8lbHJuRGhZpEF89b6xiXbeY4dSCrzM4kpDQT0UP57CdlIfEkqQSH0q5/8ceZlnygW
f9erdPmLXclbBCWdO20KPGhwcRTIPo47DZG1jUbdSk6ex6xNfCYP6GBAL2t2ew/5IlcOAtSIMIfr
BdjzVz3MtBJAcAj76n1qFtTqpZ6PayUFPiO8fiJAvA/gQYMXH7KFMibBOkDBggh5v5NUe55FEkvA
CqbgVLhpzXifepJGCYBm3veZ8E1vvzMobjYEdw65RTdi3UQArRg+X/mYwd0j6fiU6n6Yc69wZtjw
WyS/SsCkOw/gYt1xeGikzxnpZsrK/TsrFmrrd50zX2gv66ogBT9mYlA6n0pOtQQS6S2VuwtfwGoZ
mDXSJU/7gNlMjflIGZkUbWqN3WvNXmdFuLHVFcHI/0TR6uM8ehNoXgACeuqyugPxO34hnzLZKD+c
xVAgI4GKRaT+qf26UZ4ckMR7Lc36mXhwiLqU28g6aUL2CcM+CHHNDOsVC6IWj189PWMu2qxU3nPa
TsIF8YXeGkljaOmV6QOcnfETwBgaB4YUgw4nIVFgaTXrurCL9Unak9QWtf8M4c81vlZoRwjl699n
fzVF2sxhS/MgYarzrOWD0hSiljtX3+M7zsWiR5yudNl/JurY0G7ugIjlNQOFdSWeloh3oZ2gSv2e
z/5P1Yu5YPEEOKrWhkDBd7PP3sOo5dwWV//ITLZ/cgRwR2SLt+oUKCbKHJ9Seq0bVAsYr9tvcP1F
PsnGMH0wN2xkZE6/03iylhq3ZHol9uw31TuPMWRYxvKNTlSyAMbYNJ6U/9JY9N+d2pQl8ZhGY499
/EYQ1NR6PL5eJJopgE+buxVMx681Pvsj7+mgJtrrr0y9668kyC0oGSKxmdorwnyXGnRGuYS2yuXg
yk3DFc8WUMeIH0FW1DYe7ZBdi7mqQMmQNZQa1mWXmK5i7wbkq7KLjZQexqxlzVwYg8MW4u+vjtrb
vnTRGwMn7blqksvfD0ojuCSlBNRJXRZtftzgAyz5BIlckBAaNMozmcxD/Cz6xIrgST6cwGA7lPkb
J49Ak9BhI+j83jM9peu/tzbwFVdP6ytFBnuwz5KNQnr7h14SPK9nJO9ZgTTvUx50CcbT3z7PYT2/
YmU6odnrpbg0z283yhPq/xjjwAaV1wrtKDchoxpOfB4roltucjMXCFmBl/CHR4DzwN+b2iHOTAgv
Yg1qOZQ3wID85s9C0Pe0TzUN7FS9exM5scxjgMMQgGtvWssK1OHaOl8hWbMmHZPgKNWYXHTxic22
gpeI4TKpkgM9ReD8FBJ06wHID8cg17nzkXoAMNFWc23QUCOQFedY8hT2rhf7Uyx2+qbeVgG04o06
Qf8WffQ/aAQsM7neKiSkVamiG7UfOiu1byByLOtjtyxdIpP0j+2EF30XIYRg6B+8b4iTRrgoY2Sc
IhwaCyjZAVXOPOkcX4x6aAKhuN2SviAuNnDUe7cz6tXvhcfMnGIbB4C/g32mnCb7fnis7MiInjCt
vEc2AHlmL1RGY+azm3EJ2DMhXy6WKQ9+5o45B5y/VdGJE39ItlLfqDvBv7ZPBNwTGzGDhcpMa1n1
hu0NQJEHcnnCctzSMxGJnU50dQwaa6JRBrtGkL/DbDwtBR9yc0T9tuT11voBkmTEJcG/LV/y5+/b
ySAw3vRvzcUBQxDWXPPn3oS8cKosBzTituChFIS6C+Ea1AgVEgIB3VAlWEpKoCtM0tq4IJZqynqg
leYhM9Oqs26Dwwzqto9QZM+I0ScivFS/lwghzwH5GXm0/J5LqYuFkOjMyJfxpvPct6Svdo0RVvBX
RSx6mLYWv12h1L+Fx+aP70FadOMQfrTctckXkDYWGFc7AmQ6JMqNpcGTW3cUxOwE43GzdydpNTFe
Gvm46nSL0sAd8HrGFyPJWc5RpCBK0YBf3GZW2JjwQYnDsNGa7u0ePVJY1Cw3Xu5SL9p6hHAk8p7+
LKyICuq9eN5Ja6OKopOlQeX+MhnatVAV5s6BlObNuNiQFchp1oXOfGQCCm78cbFatOebaDLK7u2o
FPzx8EOy40tVlGD4jLpv+npyCJ8Gv3Xc0qKjQhipt41/yMrgm3RrI/jykMgzt7f19KmER+1qcFQp
X8CxUnnUkdE1OnbAGPiuIKx8ROIjHHtYc88tBCKVaSoweQJ7CgDI1cR013Gh0hADOKy9oQpzl0PK
FttSkvkeBgt6MRqpDYNa9OWZEloLYNKozVKm0sXaNonzszK/XsFzLFIztMIplaLCbUNdhYG3utKO
+szfS7e1Arx1SGS5tLxOaptcdl8WSO4cSPo13WVGezdH2HDhef/j4bCnWu+SpI/TB4a1/76Ef3EF
uHLdBpfvUqpcvfgc5Ve1b0zGyqk3dafnO56M4lFXYwEZ96ur1VZOIQ57A66tI/jHtlj9TIUflhAp
+wDygGrlf6ohl7w8cFJ5uv481TMuee4CU5TPyfd1xacjGOg8hpM/xx4Fb9jxYofdImeWrZWIaokn
YJtC1HZprlBJqqYYt6zJgonp2BcI4HM/jEeGLLL9OPli5k9PNLk56cjgMowF0+CI1qt5vliuTTjX
WgaYPZJMuFDdCI5E3y2bFC3yNJqKtj5Oqgf5iYB/vV9v0zmy9kAfLmMoZNG0XeKALVIHFXix6kdp
w1eom+yTE/VnZSiolhrSi+890gmgNitWz6JJThX63nuBkinaqDfSYoRZk/7IBlA2CW9VzeosgtBA
pkZrwL871Jz9m+qWEIz8B50IaIJ03cVY2CC6qNSncwZabXH22GmD6j9GQosvdMikwNojOgoaHVMw
VEpw/kD61FZz7xgxJi8JtidDK80aWMFqgB7N8iXCUlZcAKQ4jjmh/Wwip5C7L6JU6vRWScWT01og
GRJOGdsdjW8iezQxE2V9pCmVIsl18xyRvCB2Zs9aNK5RA7AGqpTA+d+y4Z0YBM30/A8w3rgq4p9N
NGQh2rj/7kOUs8+kqpXYpG4+NuJNn8Ipx1V8zBNgU0Qv89Ug8xSQIcy+Uhp2XXeJm4Z/v+7CDRsA
/zn9twWTj8b4jFqbLuKQ6ShMJdtJoIwydREu3hfX5FYsXKJlku6U9TDETQmvZ3E1u2uVQisyrHoA
RyBhDedkbagbcJUH4FYLHnsns8JbzMa+ww0faCGfTbSUSLcukjumjXAsvWqvv0egQzTRhFUEaoJc
UFR0c/q5AQXFKjB//C7toK+EGFkqKEkQxEq5fMhfBd2qyXne6+nytEstCezXKOojTzY/rNckFhYu
Qkw6PgnRjAiAQJOYhP3Kyc23f7b3/5XP2pom9SJGI+2YHLWOg+qrAbaicrWjKPanUjqmLIN7w+6w
Rmb6rD8acNjon90rOIov4IjVJV7aQUnTCF5LqCKXmtHWRzMruD+uQGvDlrB4sFw8pXr/A1WrIFzA
HbbLiC9YqE5WShp9wh9zBKy+bghtj64xwdy7p0brCH7NQ6hPs38XhTB4rOVOrWfvo5RXsE5W349X
Dbu+IzBAuWRYHMheRXNxPQMiBH9VoYbaaUdWuBpzjfVoSrnFXIZkGOohQ27bmqiTB0Xg6AVTTJLy
GEiDNDy9XZ3He3hQ259xJrOkeQNIiZl746vWXwjqKRrQldxIlkUM+aGpWHvek/9uMCiVjgdBUNV0
0wBWwLBqUtJDjznIplKfLdx2K2E75cHbL410YDHiUKeuQLRfiM73QtRVb+DIT9ax3lJD3hikWdDW
OOHmQ45Za3PkI3ZgoZ1lTVf/LWyuWLXB7WRl5hQykXdmloktDNOC0TvFZJugvWld5T2TnEJswwLU
ktLNfCZKQM+t/9MAsP4FyE4J8djvXu5z1PcNXED8qwMgTXNU9Eb6zXu2QYgUVrlI2tpWNqpFKBrm
wIgbA/jqE40RDrKb7ZPBhy+BO14e5g/1AdeB6vyVc1c6keTQdZJd09BszwIc6zHo9F0NxbJb9GaL
RPWdWCHd3y8GiN7Hnh0LEN0iBe7QRL+wf409OvfWdjD2tLiMcEOcg+phX/ToCUBywHwNVZ+fYKPf
6nuoj/tp0OOBfyKi9bg8XmzBSsfx/1uSJBnxJsjgfGzFrAYAWJPsEtz95vEZKb+WSdFPKvmY9ZJg
CkZOL6CColK8swaL3CXgM7mZ+Wf8aTDl+OqnPbYOlEPHETqpsQDd9GPcKICyknU9EpBvBip4D4Cq
FhDIajoh+WuI9gbtuTu8bDWy8DLLyRoEyx8MXeUIcdKdEg0dlSo1aA58k4FQkvhuNyQGHXMZph/T
gy4rkP/ZcEPNvZWEn9OtsWtHw0uyIBcEVDZjUASxVw+iNn6dZrJKyjSJjVZN67Zv+e4RWLrsevUN
UbWqV+dIiy4OLvVMaWXl24WS1j3Y3+CJd+R2kqTgwFWyTZpqp1ETtVxD+QVeDr7lH4tKr9XZhRRE
dTrTzCZPFmcU4UfNvRcdKwuXV+hx+UUBGYHu0U/GMnOZBAKTl0djPzlUDtP+hMJDy7Oly89SFOYq
BiLzpoG+z1pYUvUENP4SUIUS94Zho5+z2XdXCNPrHIWuh2wNNZHRRAfu1dPC5qJ3Oggd4ldUSac1
TLQ5/KX0ThbYiFS+TMU7DcFZo/fVzgIexry6+bdZ8P2lG0ShD6owXUQQI1ROfUeYu0FrtWHxe/gV
NG1tlJSWrsizEDCs9rMAZUqkrEVN4hEFT4tVpIOznIqEfuohI8huXRs9Nek+71/fGv1iFAs9Z2Sm
ThV66eMHS7P3TR9FcWFgfv7zc1ryeHR6ejb1H9ACFVXm0msfmAn9SzccqECtOkq7QfggaSORLjE5
V4WkBPsUqNK+n1j/EKmJslo5xLla3Cl4H08dCLfeydkd93saIsL2JZZSc0XRF7fRWPpfHzCPCAuE
XeXUvrt4Y1Z+rRvu50d7ndIq2YEljQlPk7JXBf1LPqkhTKRZ/3SlNYZxoj4E3kUkT/Smodxq9u91
meEEJ9KrGx/bRFOrE+jRekuGXkN6ezNncix1voZfCzEJ3wsYd5H+CTMs5Z8ALlkQ+KioKhofT1UP
+YES8cUpblGTRe0LEk4SdZv+W8CcQ+xp//bcjxL/kW4RDCLeJqLUeegQ0X2coQl2lO6XK7f+map1
FKl+vFc+w8JbCLLcW2XvuUDGiGNeuhnFQFNDK0IapS07LNC7Dw0uECox+jY+GpQ+0rSj2qZvwPwu
GU4OBI9Zhd2uQqbGzMQfyEccPX8YCD8w+pJNqIBJxBrmvkKFMXefzQ5EdzWWx1VKhRQgi/X4lAwm
Y1bS2yBHwr4W5kGRy48cGvsowIdbgGwRJwc4wFMQYeBIBCWc2hzAJy2nQGnyzoFTBKgniI3BE1dA
kx1bFXkFiWP7XqzlmyRfUObY+iT0WlHOyuecx0wTKjVl63PCo29ZVdPyljJjg//Zx30dkXzXmXE+
h/h1OYImbM1d2aRrKb5u5UUhEzWNlhvH10OleqVj4/H+Vewjc/yclZUy/fBpOXOoThzVia59foQ2
eVnp+Ut3JXUmf8G0DO8FNTdl9gTbkWqf9KOfsHfFzztzGed6FHRm1V1aCOPDdKyLzqK9g36nhYiC
1fZTyk6DxWOahUnvE0hwz6lGHpP2w6IBxyd8lYp2fr+Ucru7XXMQnUzIV1kvZLR1RFMOdjZ7TGqo
yXMDXjTQKZKBTgF8cEs7auQ37l14zBzM5p6m6+QYseQgP/jwlgVU3/4SK8nE2le48Zc2IkHZLHZa
EXoYFRjgY+TISDqapzAhhfiYeg/0lwUiAO2tqxJbJpPM1CzCzYo9be94RTYyUXxkw6EudIOvH6KR
Cw/WXo9dFq2F2D6m+f0X5WY9CQRCkI0jfPLBV3vaii1ofAuxxStovUlwVtNbhgdrW8gNN7Qo6dfD
b+1gGw0HqHEZZp/sSghVOK0onGFSUCaiITGFliWoIkXB6oPb3yaE8e6/Ng8PiAjA5eSaXTlW8AaH
0WoOUWXqxcw6a3HcuVmoHqgdhWH/QvMwOVilBetWOPsLIbacIb88MQ1CF9SwgT8TMzTYN4qMBD8L
xm8RFHwNW7UczJbsRuso78986lg+0qXxs2toc6gA9MKBeWvM5mkvJrXZMI5sBXFQ/4Ye7FIU3ebA
kz41KnbqINz7Rxh3WfersygViQS8NRzxG7Zh6xb+HaEeY1/aD2MgCH/EJw58DtHYNSv+VE4ew2GN
cIhTZEUYxeTdsveQS9ZCI+LH59dPlpds6kaNhZvoKfDc01Jq93sxAmf+Pf4Ssn66g4pzLL8m2v+A
IbLC3S4LSKxY64NjV9PPZixHo4u7AC45AzmLI/IP86ZeQpGYI+w/QcBDV3KqXE2qPRZu0NEjJBoF
btj0FA+/T5gmyk72a+Q3LFj7dpNxCEISPtA5WIrtsGE6bOYzEcFfILy3T+x0JIvjRVUjp1dTKDL5
teQt9TVjlG32SoM2rWVyuQ7dHmeIFOS194rL8itYxg0GE9pNBUIVwFk83FlhyCut0LeJiQc2eC/j
zEZ5h72aOd4XfQflEhNCosQ1KTon/LuutiiNk2L7/n/+wgKwb+pxFM3XUtzqHGYIzBtcqz9u017F
YAOS5uOV2tyArKWd+Uk6pnjB4WclkW+CpB1Tai2eyVnhlOGf4uHuTPuHC67K8W7as3praFZIw+01
PSRHi97rTWfQzLWsBsNS6vkb00xeuuqYp/C0TNoONT2UFWkCtUBePq0fg5OGMqtL4DK8xv0hhKbV
b+wRQdTpIEVdPKcYluJGc6EUISmRHBn9aGrTH9XH+T+w6K66+UHnUe73fN1TbAzSRn3P7fgKEd2A
+bNzrjKedF/M4tW+BXm/I1HP1h/953wjMO6PWt5sNJchnDiO9IaUKUJrMi2LE/UjeJWS2GnJD7W5
5ynXtA/D0+d18YSw0QyPzex4KfeEfLxbbkSi8y98as7CP+6xFuDlVYJPaGdc9CRNm6ykNpUK7jww
IdO5xLG++fNLiCRrA5+qadPX3WicGezRT2K7HR+FR3NAc54gKyGBG/2wGpqlyn09XWzzdtsiBgoc
eETu7aAIgzxEfTAAF4kSQYEbn1kK5Fq7UcgNM8Xq7OepqCo0gzBIHzsztP8giNzawjWAleMNOvGK
VosA+CF+QZY8BR1GNRHM0Th2b98ah9XHpqQbiCWMR0T/bTB65K3eaE7z+203Ff8ZPt2t52fNeqpp
ieX/FLS+FRqxFFFg+X86lzWU72mH8lYzGFEUYt/YZ/CjvklqPsX9j+Aw5fiVGrreSzM/IsHNtReV
XWT2zSzJMsTBTEcmz2kx0A5DoA/abd8fwPqeT9sbCwJaeqMPZzkSgv+BykiAEsdyvFm/nRY69yob
a1TRCy9RAg35+7ajNMD3S+A7AjrmvEU6NAiNsfoyX0Srn18ditrQ4k362d8hPWZeJvE9rxUEJ0gk
C5bbAXJzeID15vAwGgRPL3puiWAsc1IlUjdv6iGQQ5dz+rygc7gRXKJMyeHXrjYz5j0JTDJCGKNH
Y6KsrcSlLAPzjAs4GX5VcPkFxNkfYEUh8GDv+JeuRMnqg/ljgm5k57pfxB0oKkS5GT3grhN4Vjqe
fHCcAFP2FVi86Yre8ocnQ61SXMx5Vb0tr4pC3AQtW3YMVqU/05THTPhELDiIqETy+Rh9bG96NH7c
K/zKkIwI0KvTdUE0A1au1/vFaUt8g4UWSl90XXUZ8irmkWkewbAQ4//3WrIIZU9F4IxGJq11u+9L
uhL/9lcfEGjKv4lWer29RD93quh4dS4JkNHC0pDOkAVyImYGqHjyC8ZhL3u75IENRqhEyq5frk+U
v3aM9wGOMBUiJMYeyc59AcD/m+jPcMi/pWqT3mi3c0nSbJehzh8ImB7OPBAu4cCoWiviYSUFvfif
WrK1XcHYxDhZMHubZ0eSkX4hh6vVc4sxgfa7dSk1mF2n8WnzhhvhjMyNV9VRuS9bbovWe+BbEfna
gIjDQth3a6piA0okHDW8r7A97kZmMwYa9Zyk07hnRJL2BTSxo3Gdt7QP8wFgTFUegTrgWJulnrzq
Mz4NQ3WaLcha7x7ovPZOnmLeBoIM5W/frRYLFshg3au1nEW/wVtOC+E09Npd7qo3/RG37H4sJ9JK
T3AvDEQn31QVc67lTFPZDIPVrxoEZ5qBJyzt3cNdXOmlPObCI0y3fQyLjGjoi4ALhjyeyEofPiQ/
YWK9jKrTwZuImA6DpqozFQ+xkMlwORKU+ZB1I1Ma/ULjaFlNg1gf1MJzKNur/rYjOBFASvjaV1i3
E7WhpfFQ+UuhCVuFaRKq/QS4PbU8Ptu59dAJaM/XQotBZMebKniTxuQ4e9MIVMlkQSrwMSfTxW+K
w02DqkVlkpVFoHCyzRwcZn8wovrCS0WdKFocrop5Xtir7SI+DxmKePJh42OYFfJqHY6urSOKyI+l
TGWv+voTer04mStPIPdLClvXlBVgnP9qNtg6RpcM65lU1mhYliczycvK1EkNYKCp3v4E8xuStcoi
g1INZJZRAn71z9xzqft5MPCzIEuw6MkluHXxY/Rb5yBly0LjzKoTu+JGCV4rJOwjotcpY3MFvbxz
ESUGWtH9p2lrNlC/R5cIK/1S1+RUrfSKuUpY/ymxSFABMko5TkPbxWDOGGo2fNDxkutp5Hc9NgZy
KKVwaJGIWVWlT47jcLOmikAeMQZOW1KkK0Hkn7RxLD72IFody0LaZi/7/OCwphd6N3QIqFUZjMNt
cDyk3Y726wwO2AT0F47Uswytsu1FYHvycuhvLWUMRzohTaTW8xNjX4Km6ehLEGrUkmLJXS3wW2cm
SQJ2FzRr5q1SkeIjq6DIk6S3ksw1fgYp57Ct9H6gzln8zJM3Zv//NjvuECQecr1NyAlXmsJ8/fdH
VnZIiOlJ1n1V5SbCkUfFumeZIw9cQ8JN/1hi7wHapfB2ySjC5YtCJEhTxnhjUvIsKh69hAggNM2g
HFv+ApABqyJkv8LmOU5JWf0AJ3L6yv5wCvu1OWr36L2i7iTnoK+s6pGTho4CvS5rvjeLWnpHibi8
9O1nq7tpTT0TTRMR/rH3C9ECfzP4oA+rBX3PA3pQbxTXUeZ14gLPaW0paOOMH4UFrr+07H6GsCcx
r78/DcQYYw6Dk0Fgvq5PCwo2Tg0MVVKEz2L6HeuGkE5owldKzdxugIqpoQ66tNUK+y5V6y5Gw1aA
0srQVEz73Y0tImLzhPa3tZNQNamO5N8H/PJMFgUC1n0w+XS5N2UkNpPkeXMkvXlStPqZmn0f4Ase
pli0fjPrg+cXoQkaOKzGfQeX7CV8UVIEE7iu6Lk4OV130BolzxieSp+wS309bqxJb4mAIYrRCCzl
Jdam0q5gbtBCj1qSkuAK9qsaORGkvSkRdseG+nhdYkTPk0l56B570ujAVphpK5Jm9wujEixEG9Qo
keh5pXShJRw1LDGk0hx8mOr/oAdtbH4UndXT5gNSvosu0Vx59ym7uDsHe+jgxEJ3cMemFhFfRm8Y
dwz1Ujvl6kjVzMhzF9ix6NywmzMcEit3cXb3zc9YOcss0WZpU3t+s2A4PlosSTjz34AMtDFgnbuw
IiGj6fibqCf/3mQ1ZhlBhh6RPVKog+6ZaNgczWL5SUBf9CLgkm/dac94Q5SICX+QT9VSbDumxP0g
E9UeQWHqyoyojAcfWWXh/sojQxIBseJCVs++wmaL+czxosQG2iCid2Q2n5SbJVofJMMthjy1K0nd
qQ1J4g8X5DqGV3ftM7CQCKu50tx1P4rEj6/S3isj6EUX89l3+dRDqc7u+V+ISMUbgNTlxJz/0qDA
ysyeCnw3pawuDPc7bWC5Z/XHFiSbyMjQBaJPZIPsL9EfTmTHSec7odozt/ZsNu9rdj0QCuORpsQr
sd/KtHW8aOGx3ODN08BqaUKpYh1UN3l2eJN+GIOhFO8M1McXOR6wB+ysaI/Idh7SktvKOd5g0OjF
d0A2m+ajWBdrmqcmWAM/sNHJDLSRNKcfaTWdVj6hFgdjyPB/kDCLTV15gmecY0UrknET6qZgrdnm
spTtSP+M5sa5WrfvI8hLb57p9NyiITnQJSCEEBgMYO5pFh8Rk6lQAzvA3WplYCbdZpTSisuX6/ez
V5dzx0z2nELOvPHG854sH9P5hoaA1x+N3nj+l8W4VhjnxEhNM7kXHOFLst6EBO6MMyw+wH3qKodP
TBN2G78Paee/zWiRG1+EORviN3OFZgNa6qG0yS3R1KXI5JycIC+2OlzpYtWBH4qDHJj6ccfA2HHj
yiObDnDjPS/t3BIel2OmSvGdB3wX3a6J0/M6UkPcYXzyzIDY9ovel1DEpKLLTOJCCYYQfrRzppXj
1rRornrzGN48xccoiTYWl54bsDhrqMzto8GYMi41mr5hdrxyC14+6VTP7Etdtj1oZ8+wft7A/jbS
azeBjiOyR8XywiApmdlenKPLOnjy/ZpJuntopjKkE7Wx/Ht8NK9zSUt23wgqTB1rG8+CJnqMwoUO
6N9Cqj9R4vtM2+M0pGeSMJmhJCvE/ITt70SyvpUqlH2so5zPWu/1DFuLJ6JpbFFK7LkTjLVU3pYF
LYFHLcTQ2iQ7TCtXkm7i+r1jcyNDOxAbRWLEtxw4UQlo3kI5g/Nj0VJu3GXxgg2OtO3pW4PD0JqI
o9tRocgHWMhucLReUPQj8zjAAvuWOl+2G6utJCus/5iGsPRf9NA4Ie+60nYyUT09QN8H8LtSYIHX
Vlr9jCC5pPKVY5i0q+Dtcd8JfzKd1I2Tnidcd91OLSax9ju3YeEQW+8nahJEYLhLYupCCIk5e6CA
OGKLFfjhSvEy8FMp17GypolAGu+ztQE7uHRExupxZkAu5xxDlA2z+bak6BTJGSWXRu9Pd6qS/A65
4GsaXmKAwn5TsM0LSBJrpVwxxchyer9psa60jRXGacQR/TIeY2DBjZmIRaEwzHXEkf9exzNeamHL
Lttnoc6ZeSVmEGSzIZixjlaHEGmuGO8zyujEcsGNboXNv/PJ9pt66Xbrx4oMskcAqrm82G+Vf9UO
PU85+NyS6MHDKhrbF1+06J51wQ2XG9lo+uWalXhiF9vSr8XSrSN0m5UPVQEn5ZNtbSytdOsgKqhI
xtzfIqU5MQX3xNGGSrC3cqg2o8fozbyjWeT9eTIFRXbb+pRhlH2s2G3HyYVMzD9wQyKhW6iMctot
9rTrFzrZSJdjPnWzmcmX1jtMtalILD3uVJcCfQnETTBHogpe5Al5RnR+6sRDkDTwqbN7DT2Pdzdf
n2GwiSBnYWqNx8beSMxLghmW3GM+/l2awJzzILdXldl+s6HZF1hxjOHzpNPJiU1zlHA1jtidSIzS
ndP31jNPcRpWXU4lSkod/SYLFQr/64iLR++Mh2PgRTLXRIeYovq3YhMznJS9fgS0DceD2VZ6qCFD
00LClpfHTXWPUYrr88M6vh0kCuMRlCZxUBrguB8Ld7YTfDfSk3KnXt7knaQZ2c9iCYaiSZab52Va
naXCQDcXWlY+fqwi3e2Iaypl5Vmog3lHxTJbPoE34ZofbT4hv63GqAmYonuLq+o/wk3ZV4BQa8AY
A2TOXk7rR4LnI0E11BY839H4C3FuKsizhA9V6WuNZ3W69SSWmlluxyoEHTYH/75m5Q9XIJZEb1Rc
MjUrteyukswfJsgrgE0SzTvd1PQMc2Q52qdGg6/uP6Fd3GulOJd01mcaAVUunwatNxcuLCktAOdN
ZS5lAnAn7st41ruALAbR45cFFYG360PA+6Q025MSrzsg+X1mD2GH29wKHNhOxfs5XduTOoBdbHR5
R2LQ+H59IvpMK1RUHe7tpM4fhf8vomT2RArsFkyB9Elwy60hTSy6ZXEGWfsIDys5UdsOWpx/wsXf
pKu7p/sbLE3TxcKlTIJJeN15cHhrZ+cLaE1dXJ3tSdDhHYcrR6EQ8MfCuqnMtjUXRoPlohZjwiMH
0KoQ7aiGc4PsbtoZ2d3fliGsCXWjSPNIM+B32VA/hAZOHDsIRbJjjYYg1tY28VfXZ1o2IroPTkT/
/ydsgG3N7htiEI0CtZ8fmuzb9vv/5GrI+nkd1WxYuO1/P2ARR+wnYlVKjpoPJ3JXbqhP4sktPa5W
YYxfyHQEQnVDx+AWAuQypC2Eh0reGMa/HjwvxAwzSn3zBhZ/WVL5gEIVoLcQ9mzYa7Oqy5pEXc61
4br+pZk3C2nnBejHF4M/At0f0ScikQ1c8iPEyFiqQT7J3l7+0FeCJfGlLv4X00E7r2psOTTYProo
HqvI3SboMUW7SGu43YsHMu9+NDMOmv5B4/67bSvnNcc6qOpVO4//OrKBa8X/yfUYAkF3zh+viyY9
8c+dfLpbvy4BazuvSb/L67Bklet/bAqtWytZjL1YPOP22isdP6vcdbLWdfmc/2dYp7UAedVXTgNF
rwP0LYA4RkF3rljKcYKMjOJy/vi4+m5huetQ3Z8IaEKnKAsSO6IPwQ3JsGIdMABQKLIwp2Q64UIH
kPFS0x3s7nkYXXZTDvLFa+01ymxI1uyBnFyplLsdCG66LYH0kIX5ejIY5bJIrwVoVT1AJaU2L1dj
zV4P9H6Jk+oWDjy5+waqt7lYY4A7mfpnS8ttBBZSp1Ul1IzexCgvJo6DQYNLklL+wfcmf1ursa/9
yttYLmU7ZgqcsvmQwpHPDY4a4Zsk1aL0Hr9XkOArnSwF632SzzxOutePacPc2R/gY6koowA+CRA7
sNKTX6R+GhOUeaaxVr6ttfZuBKZea6jF2Ll9NPZ1zZ5tXKjTAGYdbHg34MK6q4ZQqSwaUttxS0Ae
gStr88cELZh3di1YlRLA8+mogHwcEGO9GTZXPX6TotY0178mH2UWicKmhnPODIU9PDS8Ilvaz55n
R7FiOQ6hUG/DPYYh7Z2/z7PfxC0F7YDlHAjdEB+gqkUGLnLvxt/1Xu4X0pzy+WDdH7dG7o4c6azg
y1IlOToiWiBmQJQCnQVDJYGvdnqH6jxch6Fw4P8ycTY0l6iSMg6LiUuPgU0BV7d0C/ggILJOTOrA
QOiK48AR/ez3QoLGPp5Cg+TvCPI2eS2PiY1miwQQrr5ukMYjnmhjtBPDeHHQiWc4+27SUWIHDsQN
gdxCecssvrHd5bIApwCB9C8kJXVY1X74clwKS9nCsWBbot58JFwiOOW84vZkR4ylGanu9z29BzNq
9qYFBsE42tDVt72JIVgr9p2l3/p5hnCbw1YG1vumKUD16e1CGe35cA63XCUh+8WRR/qFByzq99+H
W1yZqbU3+a5GG+CnZv8ps0xHZ0JULZYbSDDu69r2VFK3NJ2qIy+tHajHF80wi/nqxbIpz7GeqDSU
7gX5ibj95m+cXNa7IvCeSnTRKUllIvTSYuEh8vKKWqypx+oPD75Ypq/4ood9FmyD2fq0eBGfOTrc
ZNgF70UM21+4Ad9LkgjIHdAmPH7s/fk63o9PYYR46Pz0bqb7viNXZHd/vMORoOAeHchup4I/gxuE
i0GYqJghE02GOSmlCEFPAiH+xKUhOA/EoGse1Iysxmkcq5oMP88+CJ22Gv5X+BzmKryqYt9FMZEn
YqeUstWbGsJfq4fRZtL2ql/Y/TjZnfniQej7LS9om2YaL0XhmKHOtPHj20xug5lp/qPa7p8YWXLY
xNWKm6BViyZERmF15qFo4IRHBCwW0tr6yU9swt9IgfsWWP8M8tfUwMe31OgLDK4a7xBSW53ildxs
aX+Wr1PLakdKxPePLKxPnWj1kMDLyGHNgfjQGfq5B9oDc+STbhSDAtIUAGFw8abeEmRnnrhqRyNk
1lytUCK4yW2abSJJyISLQkjLJX/p+1+a7f+Vj8T081CK2oxyB/gtTHDHW6/aDrINCcYt5mzjMDsi
HHALg5jQZ02YjYmIyqYaQFxIJCrzl2nTfvh4AH/XhLA516BDgPPd75A58vpK00haWZQHkV2f47u1
247MFggBHXqX6S3Rx6kpAzzHCq5fHMejzYZ0ki7nSeM4/+4ryxKDNAWOzUpVCNFLBMZu1qDYGTJL
GxxBhdKpDUMYW8T9A3aOZ/VRKPFBd2i2qupH60NqRV35bVwGDYMckxWKsGBGmyJCAa+FovUWXAoX
jnu915TP61eeS6bN64kwdba8zbYVVXvx8r4hFAY7m+587qkJFy8NIblvgqFLwONNeFivbCGIUFVf
YCEkU6/KiI+ypHsGW6pa7zLGiuxwQWJI4ZWDBPT1iGCYHDGIaMhXP6T/Hd4jc+A6SdADLjqVeBXk
ydfw1aLJrJi/Kpbe67HOsW6sxsUoMFwxinimaW70LnED5lw2rlBRFLOzj3sv5FNsUU4jHN6zJs6j
eKoZeIOFPTs+oKnegRnR25fMri3B57Jfbfm1TQn2jNm+iCjQ2uglv/JspHmcFGGcb8NSlx27P3oG
5hP2g4NpJ3YOgIf8HWHMyrtkte6e7btFUoe7LEi+XTymABzctR410JcMN19fmPKRQo6rDA2YDDTw
UY17kbj1be05jWE1sRLXIDvHPmotKAf1/PYuD+O5e48lpt36HNDo5mnkRUHAPEMIPHuJeT4oopbS
qMkQGwcirHfwSJkC5S1QAhwMoMA+DhMDAuNU7RFtisoHWg3FuuE1q9Bvb5dCOAsqsEKmnPMWiqqW
mXOXys6qMoNwTyS6qxQOidxdkb1wSWDk0tHEB30z8c+Ll1NbdYibVYb2SppBUdupEb8Byee7f+8V
dRc6mJM3vETDlymAR6HFwXwmWngvvJoIw+khpbs2T25bOMpp7zfsrscA7mVdfxS+tXVY+yqMvUff
6ZJ+su1IEeJV1mgR4mO8Xw+K4mzBR4wli0yKbW0dGaO4z8oCeLadKMlHNvSNEsnyQqfwirjbcQFB
RSNIalgVhB1a8QFDE8tZ18ry1ymGIG0QppWSWzTaqUEdAUrKyWOsUbI387EWhSB9j011GEx/O03z
DZ7PNQH3QVwMuo/QQYEUJiZ7T+RX+JhazDANtyjAjF/8EcBOVBWfQkagKweEQKu/CYeSqxxIYPUQ
iqQGqt/QHbjwK6GuL/6qItk5uCHK4gp1CKXR3Kmo2i3JhZcFiJnT6T3RIu73OKRrFeHzxKeX5leI
Mlh6q+S9hKs4Bd8vxzrws7BUN2TQSva6qSrIu2irgGpYB0LwSotXfrd45GiOw3rHI24gyE+SUdEb
FD70RR54fICn9kwh9lvorY0JOWsNP7ZSKfGiO1OveAWSvjNUaFaxJbC1x6hEUUQ+7HXkufTFtexl
AY5m6KSZSm+70Q6AwYQ1Vc3pJfaUI+7fb8LFG7NorioK2BE1ZSRA4TGV/BB9L4qikZ+O4t53iurq
8R+Rv+JNZBoFT+7hmGVqvX5KU9Jhgu8/k12dpB8mC+Ssxon6n1lxmcISrlkGKvYut5ovNgh4v5gy
k8v5zRxzyFNiNiYIZrPp4MELxYyfH176pFjcyPm5UE3QaPzdEn4/Fas5GYIxo+nl+JDznBfdm5/p
nnlbNBiQP0QIL3ahuQsf7XL+sX+NLK+5SW3HrQb8fW8GUfYleezv3nm+UOITbuwfgCQxmoUUvGwv
JncFwbH9uBzQz5qzKMktohTQH4Hd4VKaQ0hTXtpDOnBCxPKZoBedBTuscwcqK8fptVMvS/wTWUtv
B7Ly1bbP+xyo5f+RP8YrYloo3v5/l9mxfAhhxDkV3rIBcaLRgH+9BZtHjyLP0hbWHcmyjzx0rotu
sy7N7C4/nROAy7fKahz/xd/E3eDJQr0qe1CnQhPmHOAfFHkt7WyEyJH7DuN2UDwepJx4m2PTS9AK
FRckzH6ujBjXMsUDW4JSQJu6v0XGPBvo+jbIh2+A3xBa6x29jhJdf/buQu74zLCeTajPNutjU+eh
kWdSHaHYVYllI0+c0Z4Bqq8esARh082kTYyP9VozZaoQTHpTclPSV7WM+pRWpGTQF0BS2TU8gjGA
oBichMVwk7/lmtLVJBslDoR6u+EfLC62jv8objNztGwDFwgz362oijeKY9RhHO7R7cW0WK5f++WV
+b/oH1B9142ucagwOV6+jCFPy2C6iYfxpQMaa8/mkkkDphI1yOI3nMB1gV76Z5dpV2Ao4EV7XZZO
4v0BkgzyLOJFhtd4FqquaWMXO+sr94iyjRFlICSoEOo4Fa+Dx99dlsL9NeHADT7FQJ3DKg0DYHHq
o4JwpX0cHzGA8dkhV72YxrYmPYBKBMWkoMned1gPZTkTxPpke/2bP4Mh1IPVmZriJcmt1Env8SIo
Jt9J5bk9f8aS6bZDYuBXmsLi1FhX9jhgOS/goBB+rdBnsC38HdCiGHXzatpQggV2mzgyNcy+H/ge
LcZwANiJvhzRdF4Uv7wUdH0VTojCtdKNZoOGWboChcEekHpm15JqDy+TDBl0alqGPd+hkPjUKShK
W3V6TJhYPFuyVroY+aIOmb3HHq0G4Gtd8QUKJrJwBnn2K5UuqVYWCZRXhkZ4m4X0ndm1hJXyc1v1
8tVtUgQv688DvbiWD8R6s3NpAq2aicBFw+sBJrmf+Igl4VCMZLQyVqEhdOs3gXi/dR5a6wDLRkrs
wb1k2PupO7c+T/4Vp2TrXyz1gs9+rm+wJ71R4r3WGMD9F3mo2PyTYaiuQrclJ22rU7ebhfqLRRus
G8dB9DP4TVHtzBKEAThsBggZvTVAwcuxFLck9qJ9fGfvVUmLe2LsJxMP4hwbFnIWvCWu5JcvHfIG
9oh1y2r+VXgtkxjackQ6A15c1Cx8lIfiy0DbcMWiCsELKnW45watcokN2hb1C3QE23WPVQvu192C
ieuXPa7nyhBrc/st8YzdKTb9ecwiwDzfI/WYJYdWFHwXB+0gi2S1ShTOiFshulBXHAKFq2KgHkXR
E8rw2fTDcO4VbgSepEop5m608fFq/VL4aEqwwgy7wjWwoH1HjsFSjFbWVvfU+2SLcd4E9rcpJafQ
uvkL44FzOuliOCgnpZNOckOTMHaSHSX+FRQBlblXrCPfAb9hvlaefomEYjt1JBsCHWKyxYiyLr47
Dio42e6C6MfgjzbBe/ILk8U0tf82/thUe+ImyvKsZYIvMHU5IiWKwL8utqJ3arNAf+QFQyDcFq77
Di4fcUekWPaNWxdq4hq9QJ1YrwkLR03P1Koc8+uv6PlbyYDmpTHQK/1r7QVMvIz2E7K+rguD5BtB
GuA89Q0Uma0TGVt/rFAwtoBou13J2k69R2PXQUGgQGdJrkyHbs3nFrxTjTg3e2kFPv18LFovqDLa
eWcD+tnzH7M2jQ6WSw0Y8Ondynt08n4pP0zLTJWcuf5whUEeDlkkb9PZIQYi5z1g4SS42AGYmFDu
SghKRn/mxuxHSs3auUbGo1ixPcN3ryZ8C9xHuXFdt9uNy6n+/yNJ1NDgYjicPrvCZ+fQ07CL4Avd
c5lzGkePbqlC1gUv2r7airZNJHiyvCEnTkReSFXfL6isc8whVuUTWDwPQ1j5/6z7wAuO7xIrogLw
56TgEArf3d3Eq5PVF0pjFis1C2DuW9dC5b3jjI3KCACK6hzHaSvyIMY3W/reLHa2dCRW0uRrhpuB
g9vyC1h3Glbp9cU7fp2r20rwlRt3agQGQt4eFwkvvEg1Bf6gqlJTSAbzhe8Xt9Jxk6MXVNBmh4dP
CiOucTdwFIWneqDtVsWsZkhxGRgAArwh8uqLYuQlsypY0lRaTtVOroh81EjrW5e9cIlPQlxkEzh1
LSClG9XNvBUJj23zTxIytPx445rh76PF5dn0ZnqRhq8XgPTaSbjbsUmAL9Ju37HkLOpPwaFCdRYs
Hh8+ZGjhxz3HuZ7cKEVF/Ff9Mlo1KLeab0GdVSOhpxNzeidiwQxnydBujLmUvkTV7+FtoTSNVkmn
IYYtNUJhbZB9VG9+AY9+GKGseW7+eZ53AibqYLgpUdkHe9m2Qnl9oECGjMl97f7rQuDUTe/tpyZ6
1VXha1yg0LS3DBgwqIz+dy0gXx4MwXlPsQ8wk0pHN7D0YZ86spv0NyZZ3u3H+D4HmigaQDLHsqBd
AKZMOBP4C0iJpFHl/e0WxGTi77RVyQjUW8ikcxqR263Cyc3Naq84xM6aKi2pJDRccMWqfDTZRPrv
ErgemJIIgQ/xsyCsT9Vr0Ee6cnKDYFhtIswgxzBSuIMG7XRZxRTJtz5Utt5enNOmql4kmoQmfAXP
cNZUdOcmeCr5vq54ctRqicSikd6pcUmCIn4c1mTeaIDTQqxOKnQuDaz/hrKcI7+r57WzZ1apluIZ
Ako/ITxCTX/NlUv4gb4hC01ya3eOYF3bn04LbRFUHhu03lkk9ARRQ05GXadbIoxq2FOP473meNkV
wAbMcbV7Od+cUKuN3jL2gtHv/08TpnnpyJJPYZq9okQWlYF8Q395XHxwliKXyKD7/U0Lk65cxOIF
jHXNML5wc897WePweSXSbQ8XH+rTqIpzqaaXi54DJUz8uJhXQPFm76lCgKDq1PAmeuZmpKELYAc+
wi8Hiwk5nZUWjlYvbHMiv33Fz7vqF6zCgGPhs6ngT372QoyE1ee1kcwCRxpjz5H6l0LfWPQz5Fv0
FQzMjFQIKV6auxCLztpfBvCwQmIB2ECaZ3AZBvUc478Ml6XJsFJaE4KF99jNDQsrBWMAOxo/1Hzj
i6XHhiHC3moiD/EIGqGR5N7h/xibgNdStCHFP1HorINFThSn1mWB3o7UYWqfgPAT0ckd+d+f4uTI
bOlAL/NdaqMTWVpgdxxi+iYQk8Wqb4J5WMGIRrSEgMIA7oUbSLMawG8CuWWvITyI+vIhATS72DxZ
AxfQh46pYlNmHisaazFGdBP0ekAIBxjcWeNnwuwzCmRuRRYxbgL928e1uebGTFD+J4nbT1pX0YII
JWwIK8dnQS/WLxsgiC+zd/PMSVnlxnYXTX/ZApl41nATl/u2NzXkjiM1jjw+pHBPwBH8fv1oI8WG
hyzrIUiRTERHcIRftg55TZeLnMFmCYRsua+3s+U1sGNyx5O5scbZ4OoAueP5sY5UvnPVmD71AxXc
1B5DQLDn8y3VZ1tHLCsQKoqiPitYubxQlCekNhqMTGqJcOVNYLlOgwk9S0seSgH00JSwArYGWQ4z
UrS+IySkLYJ6ZXzy0jUWM7CKHcjGPxGnXE5kh5jRrDoYwSAOtFzKZrzCRoWCL2BCfLrDDEnFFoBB
BfhkKUEDFm+VWeog0gGz35soPW2cLXpiDdPofhkQDZvvO931gazHZjNuX5APOJdXC3ucEMEmFgf3
BNwO3emWKUNBADrG8Wp0W8u2w5u6R5AGNxuefHBV47RL/Ttb9LGQEA9qz1DKrIkvNxWWUQvJ/uPv
IwMS/5l/tWiWtvhieLyUoQ+/zBkNcQx5kXxXFpFKP9xMOUaCNZcDpOpLphi/Oa965GS0kakCZJ5P
M89CY6nbWiDgpdqEnpqV5v/Jya5Ef6y0BJ2mO/EWTaYZDEevF8w8sdM/P9hNd4TplcMsQoNDs7kJ
6AjTzUjZxLifyagfqbkc0WtjwTAV+U+yuJpvUHWd1vb5G1aVxWSawOj74OHKnqQ5mUFx78lssXlo
zpk9l5HNM423S1vs0iNb/w/+HvB5mj9SQzSP1Bo5DhlMG9LItp0OlfnNWhw+wv1xPCq+qcNYkQyr
yZwREF9Y0Lq8JoZnjONDaa6IR/mmrs+UYa3CnyyTVw3QKUtWhkr76meyG3dmL0HQc2iRLNJMBKV4
I82TIoAwwgcdTKLrIal+2Cs9jX+H0T6QV1x5iEs1oKkOnofiPBEf9D1U7u6ABPSVhJfPFSyiIXzD
E7DZ3KRw61k3RE31GRGTEMFA7/fqVXu3u/iG3LUdC6WTXgcZe53GlgmbVZnNV3ZjnoANOZ9EQ+zb
fTGhEqwqCnlbA4NYCDtCw5dSO5+3aEFhYjwuqYoemI0pFnYZY+ZsThFj5ruMGQF9t7AzCWORB4Gw
koB9pLbGTn1eTPI5Q2FRHGDPOHit1bUrUFaRimTkxwSfbYuUmqzdYZ7Roz7qAZKU/GbSaYL0GPOg
YHaHJ6cNHSZus0N4bh5Z9AX8mcizHex7PQ6Jm9RwT8H3LHxQLr2hBf1GpEyRlwT45Kd9hUbN4K9R
JhuwLEUdpbHVGsrgE3GQroMOHFb+bHTbqIXpQNH6l67f1wJrYVSAjB+QInUg7EsJA99c5u0mqGxd
hpvxQHicM+QU3zIyooHsWH8IcicA+pfQtcnC5nLGBoUFO6LG3DUiT3gFeWXXtB4TV9/EA3KRmf3c
RwuVim+6FUy5D3pqPMLoXM//APZr0rgHBbWOT6JQI03xxKFj9chB5vu3MtosP8qNiRjBSl8BGMl0
+lLoifeFvmt6OZCtHPNRw9dkKD3PmV+C3v/676VkFrNRjMWx3i8+vAGSOaW/zmA6PgBir/Mgh1Hp
JWdC7APtGfTIrybyCjNbCVXeQ/dtngNJRNl08XCy2y7vtykaPAF+pTM+AwNwBccu5j7DDHK0lunT
RqaGh8F3o6pCWP6jzzXOcwbp7OcoIKPIZS2Joo0AU/KbHe8wWgsM2GHzljdwKAk3XEuleg1p+DIN
GNiNAzfYcqwUQWzTYvFhFfz43WFTrrFX3IgblNGr6D90Gm/ycszKiUtEt+KqDuaAfmUx7/bAeJXf
UP/vmYn6RFr42lM79q1iXgvye0L1dNxnXqNahlCyQsnh4gPE7yzqMOEyWrUilYbaTembc+Uzj6o/
XQTLmIZJXIrr5byD/erjqsK7ZZjiS5UZS8glIuEzCZFnCpBmRKcHfa4cuNF0CvgV0+/o+ZdXk7Xj
gxI46JqEMKV3L4hcHHsVRqCHyk6gqdJjsBnpemyq5WZH7lJvKoFkbdv+DkTbGsijoJGCvi5yt4zB
FbN5dSYwVxbkhHUTZBBG3qDBK0syCy8VYJnT/xkYLVTCxp3ikNifV/ZXmkoaKbRZeaODZ7dtyiGM
961p5+wXpkoHRIlpZ2oMFpEd8l02wtDWt8uMxV2h54A6FjhmFnWeE0g9SsiiYipe7yBrHbCzkAkK
iKvOGsIV+YCtyVofav9PRu2zuRFQHndnPn/2pX9lOSx6MxqtRV/QYa9WaubQkwIQ47MguNrHdZv8
VgR4E+QorHV2g1WUI8pC31Yg4wd5qxuYNTkzZaoS8RXAJzln4jsgf3sJc11AP0c75YPxE+C7A8sz
+NZROIvc1mDhrqsSvA0BoVtxfhcR8+I+2VMnDb9IBqgMX5VXcJIq5BSXGTKkdQW18o/xSFUMDg/W
tnRIrTpxdVX1p5dZkB0z8/Og3T1RWs4jRxKtAiMJ/iFUcvZO1eh+mAQr1E+VzdvntBoCwr7ZiyJR
UZD8qx8V8U0VnHTN2YrzNtvqNHxyg2JLnmZA1Q5PwyFIszrlWxVoQGpyFJCW9H7P088BpA6PeAoL
6hB7CIme00Zy36bYhQF1Y8Vbj6ItdKesNq2+edtBjbOGlELt+RnJVZHvcbevjX6ZYu/AzhtKgsWk
bAuJnORc1r6SNgWYmxg/80u+77JLIFR9uroq/rs/zr1GMUj8P2StPQIWtwv+kj1AWirmjhSAV8fR
yCiAKkz1jL4dBRPxpj70EE4ms/LRV5VTjEhBtfN+lFn1FK2j+I6W5zJmvQeDitZnjlWIgb/5UbsY
cnxQRvEp5Emv3qoJoPXhWE28YwkySrUqaOVVmZr6VQjA7Ip2n30bX89fem0QfJpGhkcRqz6Eh4Nz
ItfXP5xn0/V6kUTf4jE9OHCYaBNxN8PNj+C2o4rICGn0uBWGU6onJIxS3DiRyJ80hc4Lrs7d+NJp
s/WfukrMaMxCjk2har9JH+Dg5zLJYX7LFaXIashWtlQN2SgWx3eRh/whFL66FGxPxaKpSt85CZpO
YxRKFAhMPKs46q28exzk5EF2hykMg7EmDN2kCXfZPKa20/2EtHFhf88g171/mKPIdlwTtxMZ0dyG
temqSdyrqps1ME8O/bX9ONauJDxmv5Qyv2VK6EuGpeXE/oo8cJmkwZ1hzTqs2jTNMteWGSwFpbBy
QKw/1YB79IGx0NUDHHJ6RFlz4S/qk+LtrW8C1eAbf+GKR5zlz3qUrnXRtISt0jFa3v32laPzvzck
jJ8DKulH131eZuXQ/gz3lhkpLzuGizgkI+Sz1dYxf0JUcluo4sV7V0PZAsONDapHzdtZg8G15ZMo
sfycGqbmBvpV56NTKfI4mvQZ47m1sYuM7xhiVT3srXWvgAOU+uPKoZrNZ3AKozTCg2pcfnNIaUkw
rUl7UnOTETvAvAf0YDY47EgMd+hjrAJ4j1uq2dglnuvUqKHE2Dlk828pBjoGAkfKdteKeRC8VXor
mVe8Cu7hKrVvcGFDM6HI5P6U3mmSYKKHbAw+OZUzhoQ+1BmqUOM6p78p9p54ku/j5i2kdUHrijIq
M4kZgtUQD3YSVws2cYc/Fqcq5Hf2aSt5G3dgbxJTAF5Ux9yuJxdMDzbmuGu4Pr89C85MBWA2fQGa
565YMlWY7FIXgPMfeXCrkqhfEnig/DcZf6xY8x4Fb/MsHCe9UilaZfb7ThvchKPZHu7e5rlVYUT/
5hl2msfrSIKMuN7F4VZnJ3lCL6bKFumD15Dbbh1i69+x0vfCcDsfrLfaZwh98pt/8apor2o/nY9K
kODSqS984arfDqZWM5xwF3w2b9iXOb4fQRhWCXvTxNuL/Ink+CMuF/bC9dlj9M2JHWX/nm9sTUuA
qzj+5DSpsIXswUBrNvpqbcphXmeAXRXNdh2KSe+Ryjqa5ejaCXJFwL/VA5+CQ4FNXldjzFv1HsQL
Q+dvNAQ2YymuNqEujhTeskFyWD6HnqONvES1m3Lw0qB8KZ0itkP+dDFcNQSw9d1OMr7Wl49y3oDr
BWd/Se9HkvIbS+WiEOnRU9Xm5hdLvuq8JZAXeMlGXjt1oodS/nzD9KxJAvW9ihPquuhtivxb2j9Y
13Bj/f1JZCGSTOo5ZH9ZwcLmeXZzmHFniq2whpz4ADs/wJMC5rXfcweYqRbGK+8z5Vzq/kxsgR/0
E0cMDOkxKflwocmkPQHV2UNn1to28xGqN1q5B01W4A2k/sjXXFR0aTNjht6jzE3EhHLaSEOZbNd5
Yv/oVLbmcD3+W96T13CUfUxyKcZnjoo4cEtoa0Zt6abIiNl8hlz+2x/T/zYF3PJB0kSvWNVxGHbI
5xTN6byiWHSI+2ywpeeGToVi82MIsKaEuQJPbBoof9jU2hEFNFoyBhqyvPeVaav4+83VuVVwYkpB
IODIawxIv5Cy75PPbj6z0lRhnx/3xSqb4QdHSChAMsbzRSM14lca6d6/FuhvY62W1f4ZFh7Toija
q/8FpaTn6ie4KFcu6Q2A8/KRuqAV0APn3CMNU0SLLpGuUN9tuUYExEXRDDRh4uZYgqQHYoypishj
aw1mNnw6/j+m+Lf2Uzgc6tQVkjy82TegzIYuh3pIjr465a78yMWd4INKXcgw+7dtRUKSnYpZPW0R
ZbaUYjE+aItCKHC1kW5y9vvYs2MFXA+LecGjTXVFLUJedboaVTQHKK4AmTQeG3bR9441NoBajtRL
24irjrHpE4kfLXAROY6wFM72X9NmwcJNlry8KKRVxlM32J7AOjbn1qc0cq6nVGtLx7fKIw2tKfot
BKrUgTv7mPYpThhBJB3c07HeGuQ25GQlAEG5wxkfxtrviskY5Xcb4TQDej68Ah7IqSDVhrTLOHEt
Sw7CDNWwdBkkqr3PCBaTGJ0qLxw1+S3fxUgIpn3dWHfSaxw0p6mkEQCMB7DUPxqeglRpENX4v9oU
0hYlX1cWPso5liNc0x4uDKtLoIpgLIH2nBFx6KO/ugItyYLR6TFO2KQI9LVDFlj7qz8sFlMe73HS
wkJYKUCdCCULoJse0aqu8uMyz6x2jispxmV0pnDBcGhhojrf9LR0/tuj6JkACGl/sswqrh0+7vsZ
cY50o3N6OqonCpr6XoyTEMKbY/ncZ6r+ekP824gBayZz5NJkfxv4ps0BWSWkLYDGUZUxKQzckrS1
riTe1dfpaZOyzVimBdA2xtl4+ksEJXbRvHKTACLiy0Cmc7HIUK7NeM0o0JHTa7XCcGd9xkgwdxEr
SDYv79pc7K20OWQVsVmZb8l3RP9BWJTsPFGnDbP/FsRM3446t0C8MlEU4AkC0cWPT+L6kKG5XdyP
PYMR4n5cRW8tKBq0PoVWZvagUjWNKmt5Qk0RlMgzF4D85Jz2oF/9d/Gco/W1cARGCMYXQ/iB+Xkh
35IdtmzuHnpE5iN++/bYp7Vk6Kugi91idnl/bajdjfYMWBkEX3KA2HQ7zphAw+S2EOGvuXr0eo9K
RW6q3qxmnAKPV1TrpuQ5teepvPS3+Hf/p3qLKWO0tdDEB6Y+IhN2mbpR7KCSmBeCDo58m0aU/s19
byceJWD339EpmzUvS+YVK9vhLeroMklHPKTBEib9xkrBCu/jIuFZkcDMCGGYTStD37SLEp7SDXHl
evEQqgfK+rX+TpJ1vIJHFDEyVqVaCPZpxbFB8wi8iIIyPgctyH5Z2OK7A90WSybRQ/smXXw0ZKYg
/S3cKa4W7I92KaZ8vJ85uiDoHbV9LhZgr9EWixrx9Cz8zjcHKroxkltWR7RPF8aXsnMOoOKP+qYZ
/ZdVA5NtIl1B4EvpkJjyulTDUGSG4RZTbtzZaL78p/cu/ZaFS/2wqMRit5u4iETJ1eVvzhMegoa/
NNSOUutcOkVr+OydjJyytHC9r1kTZZ1z9sEs8etgX8OktSMiV8CBn3ogto1Th+HcQC16bnMtNOse
Wq+HZnadysO9I9kV7dsk2aeMLx4frATZN1pYpRq8EN5nxo59jm+W68Nptuac4Ey83oNoVHlPSy1P
N6I8dHHXNYCc9d4NW4MUfzuRHw72GFEJr0lZAoHLJ5+34GRkTvIMlgSBcDJIId2U61jyqT91ZRBD
lmp+KQbRw/vokuAL8NmxFUDWxoUFkswTZQMmSEijjDqhfMfYrvy9LXacCf9loPw1iMPmffIasAxX
R78x2DGcz1oePXNbqZ9W/S0C720QL6oGD+4++2h/6OhycZUEygziKdZudPAh7Owd1kaG0PkW7ktz
cyRbVAtv5sCR7f9nM611AkCn/edqRbKDNjL7sPGfrCpQS7sauw7o//eZ+WFa+fL+8W0rF/l+MhIX
csCBdRbSSBAneaK04cHIcnCujJUBHqdvX55vwe2ymLlMYHeD1tOLfBEQ3+3u00q65/DHjPLqLxDv
hJNkpy3rd75yqXrpFWy7s3m8uvlL/RSMcN563wq3AkE+R/q98oyEe2M5s0ZySd3Bj1BQ1KC2w/bC
LgmIX0FMyiVd5PMbo9vn6qDU1p5VBFQVs83tuieSOmP+GJNvwrBTrRF5xsRudFw90rcjyLLbM3Cy
h/KljIKcKGUAn+dj76+TwFQ/yMOjfkzt1ejkGLWrW7yD0kZgVRxgFBCe7Wi5um90rqaTMbz+OAN3
4HW+ZGH6/fHpuymkXB+qrzcBcZVBzElMki1gCuGyd7GdQWQBHUlWxTdkE7+FW2Xv5ub4xMsZSdsH
tOuLdaZCkzej+DQs5UczyhpakNsZM0CYEo+Qv841RAQqBE/4c1OFR9Km2Onsi9XZzx7ZBCPy4e9S
O3DSbTly+0gdFp6XGabF0f87zis3F/Q83m30ha8+46QZGg0MgTuGeHLV3GR2FpRGoFrq5hAR7JmU
q9WEtPhkwUCx8jicb3LKxsqeF8UrG/laym5DR2hRdgbR3g9DNrDrXtcoRYJuZCAy4QEfdIvUHSW+
s2jFwyT7mA0YXkPJ9oEZP2G9uhLNSfFMSV/kQbDIaosuhRFBLHJyOrXgKayibLH989BZk60yPVde
r64NXFa+FmbRjWsRCKhhYF1AWGCol63vpdcgON+I6SYAPd5mbiebwBqp9oOWWA+hCAAUb5X8gEyh
+iuCZxsj9ohNZ/8R2fUOdyBuqaQdWRp+XGhzf5FRn56M8DFcyFvhISvsscvymldo8x6h2IkVw5dv
y4u99tYTmA+QaozJzGK+n9F8G9EG05KiDFT0w+im0PplvKbeZieBWPmVuZOBFww4s8RcLWD9gpCQ
ylTRiqnJiCumbOSBlQWyXO2C9kkxf74hHTIQy6tmmV6PbaPN2F2caIvPkACxmzlWPRyDQNkOns0C
TCr+E557Nc1p6X4T/kmY3Z/tUbpqbhrL8E/oTlzAhPbwhQIYOrCw8uZEx2eshldgCAQZANjCCQ9N
Cu/OSdksnUSz9Lq5J7CQqh3oZeQTll+4df/f3N/7LIndbjIN9QUQboZ3uAjryi5iO4DPIyg/6mD9
6frl/JvCSHIQnAHzubma0UlI5DDa6+YorwtqRkrSeo3RZGctuAk54dNU2Lo4ExBpXtbVrcGa+jB6
/u5ivxlnNiU7R0eoIbZhNfZP/pRLrapHz9NnHBS4AuN3+fjdGdrtA0HO9+Xt3gX1/bzVlnxS/YIy
DG05fLL+ih6lwccFRXlN25ZiiTDacURnWtMBPM4bgQdRJw+Vx7V0ZU8Nj4rj1irDY77BK9rv3Dmp
7zPgiX7gU2PtO+ltN57EMeCR9R3naQ9uPUHEh6Pkkx6eh5qDjUcaaRxBz9JCsqLFFmnOCxBk2y3G
R8V+WfPo4PUaKeeAZg+HxWHbxrR3LCANTC0Zu9aa2/FRxzf5FMc8O2xo0rRB7ejZl8OTpqmmG7AW
aApIFvWK+4HRKJGPcxM6eZaqnofChgakU/TcdJy75BsM3LIM8+F/0RpdlzXw1rmhV/oPbQQYzGz7
hn7znDhm+uCM70PgO6/C8KExb3un8sQlWR+X7cWUtbYdrAXM0NWI1zVjsHEP2BYIxoH1/U0G0p0O
V04LyVweJn4cQjvBayF4BGwk5zCnHJwRk1WZHxh17bWDF0YPWON2o9lux/Ml8i9CAOi8vW6PS57F
chSuCTC9CkjEj/hb76WdMbCGrUvFnxLOZZNhJVoJ/0mwdk5KE4A+HV+fV8Of6xGySHldt8iFfHiw
OMpMY6DHXUdGFju38ZxGOUpvpIMQnnrKEm8b/yy+/h53ckoWH3LXsE1h+oTIDeqNLphZvVDjQSkH
7z4Hjv1wMCiHVnZ7PTVpn1zDCRissdf7KpXgEjbnyCcFfqpFIp5uJFlaO/iNPsW5nshJ7snE1rJi
7EQ3+IOhh3omucVFKHCmcDcOLGGH4yduuz8i1cB8hFQz185NcQiF/vDX1EF/v5N9jawQYYJ7fzWX
Yv4hO4zO78dkv9Jt1+nq9BpiFhEBbWPZGwtzA6n5HtKv+aKybtgxl4g8p/R+PgMGNvghRMr5KRXA
ue6QHul5mPRB7rjoU3ct2xVAs8Zr/pymf0jDCqrhCKsXaM5PfxVjeVZrIhT/3cxqNBSbShRV+mtr
3vaopyZVVSbO/FvcXT/OmSA/4pyIdZ43Tp0DRRaZnw0vE8HHeEI7Kl2Hmm+/FJaCKxQxtlxjvt3C
rZ2eGdL84EPNxtPwRZJpM+2hioiqVBjxTxI4/j14a2uXinzW66hj7J2ZFPbKZAQMV6qBKY0uOcFZ
Ic6g4hZaYXcVn5MAlO1CEGMsEfHugq14xyWp9nElj1aUWbW4Q2M1zXIj79GeRwPlZ9GFzXGOabaM
mtEJAJ+YL5bdSG1cm4foSaky0YifOGXMMVLz8VO+bi2cUE1isk3X2VaVgRxJoLql8Pz2S/KoqTVI
An/J6EMvtEN+Jpco3T1q0UVbeRSL7oVEzqrxIsKVUWZuGEfAf+aWAl0CrI95vFQZyhFkfKlGqdUZ
ZDfnG5D/cAoSu34TyXUOF3OO2gZD5nHuj74X+N9YwrWAGdiELfXXQw8fTB3EkonilF6E8Kejjm80
6UWcv2/7o7Nd+5D5j5B5SXiiwWiAnekxFNP9iK6RcZGXp2mcttLx2eoKKmbSpAlRZnBGXZFabs5B
qZNrQCxUZ8yPMi3am8KxGyVkSqeQDfs5MhpHFJG4OEvVo1yZa6fIBNkvhGZbkyKdm8bYPwfHGllx
1o8hITJw7OJXdbaqGM0pTWTr67HtI3r5zBnFlQ+dw4sZObGNrymKwPbqdJ2wi+8Gws5aJTrQiDct
bU3wpLWYZf5tOccqVntZvNrseYhP1g1myZFEDrbgE9OHtLR7ocV9eWJNUIab7V86bmfpjRsRWImL
zd/eJQRRepeynGfbrUaaNyuwwF98NLJXfmO/yAX4Qmos6JY0+nm5SeOsOtM0vIMzHc+JHLtPmEC8
ycY7BagPtV+viGHYv6NQhuk8ocHfLAWv3VclWyi8KJr7l5irswzCzv6Ya2i2bjAJ26BILAXNWN2C
PgLE2h/2ghIlMrEinms+z0uYy/m9h/oBruPxCPpjcIA+N+47wDNiFz13tzGx+KQkdlwm/PS89wx0
cfTnzKujgZivU8LmkXY9G0ITuYYOw6T0MrfG5YGkG7WYTqW8cLqFj3HaNOEp9stYBmikYoj0Jhuz
yYKBIfLPTyZShJ7OC+MkUBe/rZUNuNEacQy4zx8Er/xUNshhkvRqdasEbXqfxj7BOrc/AT3ykdL8
pFB7oMKOCXWrUHHTEu0qiK3/L/7rpBOzydp8fCRcsznrqQEzAKBDPcZIX4VDL8gq8roDDZrc/uKP
dDZSof9ZIF1XEsmVw1IiOe9YEi5ZSplgCf3YR9DaDSWhyduHj+0eShK/g8ZDqEveRqaIvYK8tCzu
FRBnDoNG0ztRT0EJJbM224PLilomBjf6JeP34QUwq6oquBakIkp6v6pzZ/XUhBGZ5aqi+iGoZfb5
yI10O7UgEqA54aFcuKu2kkS0k09BZDcMAzF1lWVa2ou48YPWGThEU/mngciSDJ/432n3x4vRWRy4
GD515OtxEd+Zo52Qcb+wfL2tYdDeAon4eA/xbaH0/v2RCXNEH6sRUXg5VnH6kTtc1cchRU3kyiA0
r9HirxVoXJoTa4l77fP0SUwFC09MpjpHAgkAmQZyGm3ozhognAVTCof8KjirH9UmXIDlYYmsRrqB
E1nR8Py2fGmcCHa9yR1JiU4eaUBa0A3CJmki1eHK3WG9WxThSMo+O+pua5iZtRvlO2FP/8DOj65i
ysLvxFhFEUqPyiHjeYdXxH3KNOM8UoG+4BPMOIAH5C31bNAwDrIy9O0l/gHs3zR/F2MfgpZxe+K7
Wxyy6Um0qWizlxhT3lb15swQEMohiVUTTPoJtOha/1ohNUTMxjiZKkkq/4ErsFbEi8Rx/oDds3M2
YbpnIUUXPxo6suKsLtNBFXj8t2qw9TbZf4XBlwCCNtIupkAAeZk22T53sFZYwqaGUFpDnGHhImhs
Js56zJwtzTvm+zHfgo/ejU5kMnUBaZ1s0xsnqW3JyPhW9vkZ53NbeDOnfLgPAkzoA3ob3Vp/4NMX
vfLe77Q17Lh9L0vHcUBVj7OZURAFUbk/da0RjRa2bpFA1lzQI6ovxTcQPTMyF1dE+cQJSOWQWR0y
K+tXEMoIEupHhnzA6v3BbpK/mOK+7pwQ3XVFVxk5y/GVIfejy6Hi/5jt8oDuXq4x8WDIq4ZlnqFf
qr1SG0ffmgqy5sPjGUUhQzkndoCTMZU3pRxZVh9aJW16k403uqOKXgW+lSQogjT+zpYbL0gGJMzK
HpugoDoR1rXZfLWOGV3/4SRk5ERbK6gP5qPQygq7aGD6bzLhBofkL+ujzntahRP9a8ZWUhYLUxW3
JmLrTUp10jAguWNU2kneC/pXxG4smjPlm6KS/vpsUlZFEmkwEk3F+LANLt3CPmj10D1vOQ/M8V0Z
yp1m0zQ+7os+bN5mePW+VD6TPLFq/NFdSPV4CTRCxxspUsvdpmF7MMZp6kBU0AneVu1jyHUVGUjV
w4pAwKDG+Y92vqUvcmiRgTwqfd5Ia2m1XEZe2PJTpJDxBffiwyO+QTD96I1NgIb+9BhozZhVvzSR
LiE61onjmSGZZ/vvZAxofEbApzUuZw/32FgCGqezhGq5sFEpIIvcebUGFU+9VKjzCQsXDvxoB/Sj
p0VwpoaNzokhDHz19bcnRnRgsmk20QS7RGSs24qXOmzaczNAuabKejMz23SuD7kNLjLSy1c/8b8s
rl9Ieiy4dkKnZRYArTSbupYnsjvfe/M2V5eW5itTXyt32RoA0JURVXJ8uKMmm0PzHOzOe7z1U/wv
hLLxt/LBOHMliTslRCeGszHT8YKU6RFT+zaxXc7hOtmbcqdjuLXRc51mwbD5sHVA51+3E2DwSfNZ
H/7iUUNY2XAAYZawUtSARzLSk2ZtZFbj7h3PhzzpS12iUM6Tpshl4I9VdvCoqqb71LJFffpPC5fY
CnrTaHzrvdRs/mTDw0/A8ogqL/h1uw1k8qviCTNsOCVkuqf9F8HWRQCypiEPouf1/3VLRDAE50yf
X4NBdl6WRT5n0yhSRjyPNh9m5oWhfZwoczykUR1CJvQ2lA6UqsMHo4k8nwJH/V5LS+wn63Cw/Z+K
jmwLlunq2PEkXRYow4vgtRFgNx+YqBV8EDEKkAFsmVnMBNZMcmA0Ge0IXaVJFnN/mvwFZ0Me3HbW
7cbMvaAEbFFaZ+s4H886lWq7ZoAdTLTBmmBEbuEJoHX7gtaUlWsuSHeKFgTQHsrkDqQj87nbT30i
GhPB9qG0efwixjm5g7F0qiJPUXpAeWYf5YlAnl721mSFnK5W2ErpJ7ZJQkKyhpmOK2jo8MGFjJ6D
hnWtnm2st6i40dsRAVOQ6qyNWzgw3nWzj3BzldzfiPnF3sYksndJfe6tNj47czCUqyN+X4ShUbqq
tyHEwAe64mPmIt6Um/B9OoBlKLngOPYZ5iWmVbhCeLtuYtDRg1HJnIKZlLBcgHitaMVv8UOIErZ2
SL/MmTcTU0rN6McUYtQgJaUpTZ+pkCFN591ZUvoHGAoHkvb2yINfGSkQbWDYGkmjqHY81DA5Wtox
akfCCAA90zefkh9uaCiMtej/aqmpwQ5zw8xrwKML988VYsLSRJl2uNIggbGL9qpxUdYe6WDaqFob
zNwInxCKIKk6UhlgOJunTU6qY/GH5/bZj9nI+Gg4AWRK4NuR2/v86yruPOo90sYjk8Lvq5iEABYw
1EqLkaGTf5WH3XSWQDoNeswzpNPwuj//91Bij6u+WcZ5Q+gLx79LLwq5qdiVer2owZPGZa4VxePV
d5kN5YYE9T9Z0x2f5ejiPXeFphs/Ri9xdwM6h4goctGrg5FOIIONwRhRxoJdJAheLyO0cKjFMPQ7
ZOAHGUW1XLhbDcmE3VRX8j/reHPGkepTFtVPveQKmtUBFUJGQKR6e55yysE9L7SgD6KuRL9y0wXu
O1I50wD/eqNNd7ufkv3+hyAdDiVm18e3yXAkNgjswKDShgez6Jj4Jf+zzc3ExqpjQtBSht361ve5
hgDHHK80tS1aWayYfkOx5EMgdl95uBpjga0IWVmy0OIUxY0BvTWHUVBmrkKP9yuNmhOxE791SLu3
8T0gcLSMwNQ0Fv18L1CxHWb7k1fXABRtM4YSpmo4A2fPKpPOkuk/SLSKBQJdsBI3qaIBCl+TB1mX
ZuWK5Eyry7J/FRPJp2Cff/sOaqpiTMgbqP+FFCpzYT9IpfBMmW7Sv9ZI8numwouYJcpTtrr/gSVO
3G/adiTLLiGstIvwSR5h37b8WWZyiyEZCksuT0QjZL0PxcTRjZNJ2HYG3S1bOrqbsKEsNg3K46VK
hHVmmGY3iIgzn+9mHTJ+iK6nekk9HzVMwBybefpV1c7F9Xo+ElwsKlwdwZmrTcagn/mc5fftyfAC
gNoZPXHQO00oo5hO0JqyYBY9j5ggEiywpF5Fgxv+ddO0MU36YPhLOwSBgsV9LXMjms72U5Zxw78J
t2STSVPRjyFDKLhzR8BwBS7icyx7urWXSeAW3eww5yMTQLJHBlq02jvuTCBtKExi+PNIxk7X5Wjn
r3uhHadybUD74h3QyrSAaYNOM8HIM0b92BE5xX4ajP8fcu6YN2/CKLuhtNDuBS9mnDmLLZqwuBb8
DkVFbdDUQhaffhI+qenOMpNDcnJWLzb+/1647I3PTuLA6o2/1umhj7RCOFpJUaMxtEKJCDhWWob0
qjudTLXcRsXd+ICM/tF3XsNXwKNchbzQTzNKn42qIbbdytBUhU8UG2FJw8RIs2sM7LUku2pBSI1v
8ctJfBfQva0TfNTBkGQ8wuDx13Xsv3YeCEczgkhtFrepAhWT7RndcE1ZljXg005A67XDMzkXmSYT
pGabHxlzF1DURsDxaUxLknLiVsUECGc8UzDl+RI4x0v+ZMbqFafSikeVjmEsZIGqrwu3fpROQtGM
3kssZzWY6Vxi5NIXr3bSHiw1tPKuWgHnvjM4+kn8sW1wDR0/L5Qu0eWkyTiGRVhT56j0jgkBo3+H
ykaa1UW+hH0A5DX5Ff99FI8M/ouvxpKj+522CaYI5RBUpBB4DAzTyTVt9nCRbV4Wb38S4THESRp5
qstRfcvqiE8hUQDzTKg4LotkDsmgyW40Zoqv+sNdLBt01+uhO2H7q5V1QIhRkCIwiWCwYhvUwdgM
MJ8TlOJLBkaXssySFSxxqSoL8vNEsqsbrrH2q1Rpri8pgg+8LdDOkEN5GG+XneyafXkMOoPHZvS7
bMS8NzyGy215JK98qWErW2NoUX8UTSAl/9LSsVfiJh+kmoXeIB2g1rhJPy9jLLu6ZiJXxgM+mJQn
XhxZ8gyLDYJauEjtdomKA/rbsOCGqqPiEDVQHUosaQ7bHd5SRfQ5SUiqpgeax3t+w3gb0OiqNNPw
yhvH7U0d51amiH1l+d9LX7Fq1oYml4M7BdWgnXVD5AKiHBYTghLbn+6DQzat7BjMnz3LbofpLyTr
/Wu4X/MNzeR3pL+eQklTWEu3b6xmX/yLuElVDPnBF9oJ+BCiGtPW8utC0ah4yUrb7kccpeip9Xpb
blf2hxqegRe3w4M1Wnnm1hczYRx+S/ULO4Pll1TMnzkUTJT9sUt/Cb089X/kpOj8auif5kYs5h0s
ITQ1FCXRFmkx3EGdpfdzZu/F508wfGgT95Xrs2NXitrHvvGioTcadwEGuQJdi/8xudKseotn69sw
nRfQCG7mCU8wVz6+GGDErGp1LjbHGv3aVVH8/9+edG0UXM/Ee5GrOwuE+arcu69wgEGIYXUUU60S
PhqdfhrXBZyyBl5HP78tKHGIR5kzrNPEGleWJX/zARO+bugB2Rqh+BUetcoxvCRPT8iPiGKE+fmR
qZIruX/1fxI62UjuCEI8X7mLytn48frm3ROn4lNaZWREefII4s1T1+i9YgyCvTvM+Gdn/5jC0PET
FVuu0qezMDdu81LmDFDfV4/m+E8/IslXMUaeIDdNoh/0g6w020E/dlo1AiLjKjgAkllS7YBeWwD8
jrmNCVMWzBxea48esVArLbw2PvlBQTXb3aH0fzahj5jsoa1ElJXBH14I+qbrZJLxmopB1sJBRzZ+
Nq2Jowkzsn9a3t1VqE7hrpaL3QYKzkf/s8aEOi46a2XnhshoyPyCjAoKkX0q+NpC92mz3mcVsnXx
u/n/QwVM5rOnUj/oczIvNn6GzxKhDhLXEtVBiBzwBTVcSF2yMMncuw21crWCDAbzIjtYJkE/+C5r
HFMh6nd+wobqeW5DVRRK15eecOQzz0ZYa0s8IRqXuyV1vhfj8Xzjl0JVSqLU5PMNcMagVB/psFOV
Wecz2k2RmkOzzxKVxWQs8GCp6qIYVPjkCYwhDlmTRQbcCCOBX7PT5YPY4KAazlX1+xtU7TixKXeJ
JRlZBdji5HooNZukp4IheFJQJc/MDQyxFJGHj472gLodZWqFGvtnebtRM26nG1iimsdsekV2UjOY
8G2kUVa7WQSPZ+Y0G7SPzjnjnkFgpOIve+l8nbZZPhv+FvbDSSYeI5gQ6WNT8k/Ce24698qUHTDu
igGkJjaJzdk2TvWKtd18qY74M//Gi7z0RzHeZN45MO9EsfnsJ6LySgLvueN+6MQO8uVgzf+mA4WO
1sH4ddA35V72j6rII+oMC4HS4AfdRKP+0224oWnLl8kZyqPq/CMy5TIk9DSeAiLm8okF8gNyb3lz
TFsx0QEebxWuxprazCJFMdb2jzHBPaNRbdBB3cvQ4IVaePPtrQ2/GbdduJfON8Tqgl84tZ/WzIVG
uHoho6B8YT0kI7KWoxK1pGscF6rPSev8ubWWhuxcRTLs966J0bVENh7jCFQBk+GChLHiORY9wSmP
k7jeMFpehtAIF0jLQPrz6Hfpa29NQ/cAP2VcaEu6ZzBdIILXjUglZI38R2vB9zUEHUvTOYsNWSs2
ddQXhjeltwOV32bI/HFXK3Elwpe7u9ufOSxU43kpHotLFlpwVOrs8eOyrwq+YLVxARkkiIbrgDYH
lgXsektIDH1koWqeatnFeO5wxr35tlvYwLUOIxYJ6YjKmI6M/lpUfuhTbnY6jEOPZ5cXF9l/7BpK
SJZdOGBLjLJhCsxxhejZSjaMwsMEcsDxGoyXI6tX4fL6DadOlz3Y+rwYZVIbCVZXN2u1KQFex+q1
VPoFL3OQQHXN4veME7RRLaJgsEG1o701ZtuOHufnMZo7W3LPS+f16ymgn0C7t9LcH37HzGzBkc+f
vNO9YoB6JL6YgZLKidnmDYvYOVyyfLlq2LVC2DUZfjBNo/lkLs83nDocnvsWWFg+bzG4bi4e7gLb
93eVjhQPkL5HK4yJ9y3jWaBT6jig6P71EbrWbQ7Yud7Ub/RX6M+4ouHuDUCiCFJ6uTaDS5+apy0U
PYRJWlwVmBnU1wxhtSs1yFwOLeQoE+4gyatR9F4aNVKiRwimIH6jk9bzGgTpolPND2R7WyXFo2sC
jVhJ7OYRaJU56n6eC40QJIZwxrRFpSb1fPUn/wmDmAdsqKeNxUU9/OwmYvxZphYlwL3IWBgLdvRV
Z4CCQr9Lm9DlaOSYKqnf9ym5XYAC4o0octJS0/wsP+aiVvFLZyNUkdKR3VWxfsLywVgf1/oHxdSr
2fjhevpzr5MtLVDKY84Uevh5KqE7mttsgrtRCfc1Il0TnkyZgHLNBKzab3m3L4UAFOWpHaWYfRup
a5LE2d67Y24l+viM5g/dtf8yiEjfz+lHCFIoQzS4md2lNFVZ+eYIwRUc5AuazEpgJitdQ8Qpqdi1
Wxr37Z0pOBoClKYU528FfZWp3VvNMggC5BHNV/2HiVmBZUvH2VyuYV6x+zps5SrSfgQ/+yxsSUgM
bawV37PNPTKZhVHsinKDtRISPNjyGjb6REimC3Fil09nFZ2WhPN/LcSRvx4KHh3eGhpgliud8vY8
D0R0qBtjA7O6jsGaRKIsqjQEmUhRzkBBDhLUGUMGNDs1NYWvTS67yLqTh0T4YEYjKrmuiY6p/Kmd
tfr3cdbD80unwntz8/Z0SoBXG58BdD1/oL6G+iG2LPUb/6aIPWEEmdNxrbFL5JTduz6ZThlCQjqZ
cNRXCg9Zh7CE/sgtWe5YBfjtMEoHg+tvrkoOORA5pVL3GmJQ78OUvRcU4eqirCSEwB0xNyspE1NY
vCGGDd0AVV0m1eeSUWOzlWqUzXl5rUdNDKZi7AyvmJZ0kD6pCNjX4NMIYx8r8/zJMyOCCouwwvDZ
tzvILXwA1yLTBo6KtJ73yxoOobwNuTBb9uNTHtSWQKkJ5qZRKad6CmsmqIbf5zxDKbyQBTNf0j+L
o3SvYEOzM1mFOxDCvtyz2E8d9hlKKSbnKLLUBP6XGAaEruFxVd0cBmbyBxjeX++7GshW4YOjOjaK
+uTI0jyx0xW7RtJkyGY7zP9tiyLe55zbHit+bX1cGGwmmKR0CZ8q72KwH6Zp2NgBabXm4Yw3x+UN
oLMjFysYcxpb/nAvqqf02I7nofukyD2vbH26jvr1elpeKUEM323kX17dQ0tWEAX4enF0R/s8dDZ4
lbQnifjwNwroAtStejZN3G41WgRBDVeo/kPsv1SN77ZBitdKCP3gdjvplSz01J2lU0FRmMvkIJir
cFovN99sZGwczsmlqLbmNk4lX7eGu8s+pLrNmUlBXhSxN/0c6xpEnAXm2dQ611zQorNtgVT7nGbD
3r5Ilo/Up+zTNWpKIx/D/Flne40Ix5AiGQjreFQR0PME7KBQE3xFNlwJzCRA5UJxwOLN1ifT4azZ
fb87Y6wgpqyZoOeZy4Qr9fEyiTyaabN3UpuAatNrVGUQpa1yh2UCLO+P3CQBNcP+OaMFBA5Ici74
suwQXHjd/KeUMLd6Tv5UGid4HmgQy4l2DhTkKNOqcyf3BAzv692YzLCYRKrFEcF2j+cegKMqeflX
5oeqQ/xeydzEwpdgJMLo2OA62W8Olf610Ml7vSfsOpMvFMqNbwVbRWEDNwaVqFw4AYuI//IGJYv1
15k22R5S8YCBfrB1LAoB7vdFm5j+wyUB57n6RwFprCKR3BYa3LDqydyOBTx+sAouRj3pVDdKRbfe
6rVZ+NWL2vFEPqk27ZKjj6i09R3VvdgBE0ms9g4uotUAwgX4CIAxH5TN8Q36FwrxyoOXaXqh0udL
6f7n432cfc9yLA4pXQ2bW8yy2Ihm7jDzug+KM7/9u3SfPuItkWIHfKPGpMmxBZ8XJ5HtvtxnZwaa
zm4wGwsWzn1hQMQ0TBB7VM0dCZkWgxQTZxkFPqrsxZGgq5mEjyv5hIx4qAZbuR2FKUj/FJvOX8Z0
mlv5V6u+ckr3M++kK93R1mwIjdT2upBIDK9G+yNEBX0Ews4iTtXYBbqzBc1YUgc7D9VMeUEw6HgD
hNj+FIpzx0n3BLcATIDaeIkXIHKbs8Oqi33YN9cN5jwoRWMGYRHwnog2G6Y3e5/qg0qkC3saueeu
aEWAi3QkHAOBysjo4TOoOkBLZsq2ZIsQrw2/nrRk1BuHuostkvbAnJh6yftJJHd3/KkLjBuhwuf0
D5SB1DDwumJb7M3jANAFUqia5njTfjP80R1q3aipbGH8MXYgzwG2wvANm339J+tl1SbblxuZEqFG
HYLAbfUzCN3WSb4rlsQIzZYA6p4EyP79+lad2On0iCpolfvmms2Nl8ssMzoiLCKFi+rhLvUoJDbe
W7DWqtYoeu+WoM7M8EPBnxNb2C87vOosLrti2A2JVUiXrEui9a6sVfzPGf1Oh+NFGmMDie3ll1Dx
STd5hGqvWI67fL/tmjVtXOMyx9qaLFHOkWwB9vBNqycCeFfSsv/UEaUdoFhN2yTR8EFEOtgGs/p+
2JSM3HUJTHwYnfhEY8CaBtw/Fvz1ZFHb5/R84PjP/kDM9f02eQXSvy+DmWPTwcvF/HVb3kQKVFZF
3/plsIYYcVVhsh4trPQlFRE61UXLNeFBbFWmw5sHCwxnA7C1q0E1q7O2ZvC73DO3M6fNsYdZ6MbQ
SzNmmtJwX+Dl7EAaU0P72E67KbrUGuEtQBMH3RUSZOusn5CUA2+0wsSAOnEHSowJkChErNT5oJha
FI8q0zKuonjnJQELIOTtdzaquD9yXe36FtjNMurBNTUthntiCVi21dbzoeQzLm58x3uwr+NlI9d6
iMFLwp6sTxlHENAs2T+WkkbqFdl8+OtfP4vVwGEsm82lgY6BdbPLoGcZaFWX4l20Cw1AMq4K2dHe
qAgW90HoQn21lndxoNf+gzY6f1pjtQFE3Ds0r/venTlcos2KhWUjiMi79gmNctzphfSB5z8Ak8+h
PQx3Sw/idXGQEsmFYJq3F029Jn4YgNcksmxytnTdadFHnuqmrkUDn3L3Fahiyqdk9lgdI45RQQq7
DehjG3ceKYLDLtWdBZfbudZFUtwsfdDOtn9sckJKiovMZJQJeEpmdOh6HGt0l0zAcJkltFPmgj7q
un0dUGZLLfmCImXch0BJ3CaE0UP77MxzZdh6bCtmgcAGcMigcxDC66LnJUADw16m35YsB1ZHXU2a
kWRrUjx9iXVrJqfs/fJmOD6bNGG7yflSuquzH6uHdUIfoDJQYDxUGH/Fg/OWu86zq/Sq/yDW+7aV
acHfRlF0acpDTEwbN9Izci5r/1hl2rF9M8Wv2wE/90P+6Bwsd8LiGaOQAfH7/K1zXrkkS2uPByQo
WSU8ZTeuQTDZc5CnldDgfCkxvgoUn07W30KptlDzhM4l+JamvcrR3hsoyw+ksMfLwjD4DAFh7LpQ
nDWQPwtc03qCm+esKQ68NTnFuZt9Gd27BFEM/pO5tOC3dsXf9fEGiYDXv2Jc4mgtG/T6GUPdGOsg
v+bHQtZZHKO+NMvnZhWDYmJl39ROZ7XKfPyiv0SnO8ULEELfzFq9dJ0o8zC2R1jIJwW1YQNahftu
FE2EEfGJVUffw+AMeZFRbLstQDer6MwmChIsBxtAFLm+ULXQBU+Ch9P5Y6czPCFGMLBiChqb9Y5C
mX0O8MOVQqU9TbYlXmSwf0SZt4HdKpBLxN1XZlFrZ8MarIvslnYlJEV6qswbD0glptLlKGvEJWT0
cy/mYTy2+tBROpx/ZprOWXemzK6lQKU6QaS5NM0yt7S9j/BiF3cgEGeLrKD3H1FxUpmAcXgiwHQZ
TnnIsKXP4Vz5JCfXtagPUmt3fSxBucE2HHQIK3dRcJO9btRC51QGi5RgHUK5PRtDwyHS+7ZH+vEm
AQu5OpT60GhUYRoa5PWPt3/5x12faAIoGcsDkbXf/k4Ny7yqmoALoXqVx6r1/h6ff07jdiBPvN4j
rH/tB+q5ic+V/KP3FFBObrK9D65QWlgROJg3J/L08Kb1mzT6EN3+lT2xbW3z+PVk/P2Qn4hYwYbc
RWxQDANZxnzk7UVRchZ2y7oBS/wFWpgaKHGKeEI2vWu2Yk3zORh5F8VBWNZV0qs7Omfj8OeHuwT1
PNuFTTqARAefTEvBK4cTPYF/8itF1l/jnCChqoXnmt187qarAFX0kyDGr8nrR6JgQ2i95g1OPjnI
FDeQevnqdrZMC3OBxDU5YHsd+kKuCevi176MpfytBviey6zG+xxmtAIX28RVkqq4AWjcrrUpUMd4
w1sEKaIr4hyf4uLw3dDwhIBbd4IyNjp3Dx58DnzPWIjn1S9MJRYr7Bh4WAp4JatvIkL2ewnBNZiO
buMLBne+jZliR30LaMwkbo3H4NLSuLzRocX24YHLPeJ/JZXs1X5XxIznVoxDZ7g0p7xDUYNFe/EN
zAoZk9qnQTQxTbl0L5z7ovukwymYbOIE9JG8Uf1jpCfca+pvzYWmTssWvxBItUFR3198GIDdU+Sx
mIbaDpAkxICpbLpA8Da9Cr6995z+zR6UMiY1FB7Zl0hr5LGfxQvVt6KMW5AJXZ7oYjmiTg+UUoPP
9MKWkIHNc7QLPSCgiZpbD1D6a7BIoFEFmcVwkrKmwSJTJtEl9hJyLMkW9LLlVtjLPKws+Sr7IB6J
RZyP0F/mRPvPJ6E49mu73GcLLs29Pq8jBqMnZUgi/QXO2Br0r/x3bIyIvQ27PtrqqoWXcj1p5cJf
Cow6hlMeepZhEE/ivW4AZsK+kxYTWs/0Y0drNBj5yi3ZtDApjA2vTIUlpFynvUBqVwAwWPJ4vukS
nAbWh0gTXsU6lQOJw28ObFk9lsmL8wX67m3J9yD2VqlvIOsFt/eYYflT3SgMJbW2QT1slJsYlifL
451Pf+g6Uwo033rRvs2RkXNC+PhdW0wQ3t6k9eDe3MI1F9XcUi+EymbYN5urJE4WPp1m3To/PhHp
4BTAIbNa9GDrCag349LwRDgEiwDC3OBj5QA42m2X3D9nOVKiYGJFdNGL+Ui0/7zTNW1y2H4ybrXZ
3iLKwbpq77YRRTODRGYTruLWOTzpnGNB8MljoUltvUMDuaxHocFOldJ6gzvh2ENPHCsn+buu3r5+
ys2dD3qgJk4odTJpyEf6K7YYnPajNsWVse8wPqAPIgJBbTzXXQD7C6qY2p19BhSruFqW51DeFxaY
HjqEF25AA2KLVBtAj4bWyVTgfjEADRL3C16k3Yqh05lgzkZ5fJtbKnnaPqKO4TVi42cjRo3FerB2
J7dl3bT24boXI2KDwwsXXJ5NeaFnKsxnO+GJJ/wVO0J4hoEzCWzeVxkUQau7znYfPSE+C3dz+d1o
unXfaerRXPBDS3ou+mX4jrpORGvvEFuhkyUE5GLeUHusobd33qVWtolVbl3sG9JDSy9JR8gDNe6e
2OSDN2W9A4bkPXxNcMxilV3UrV6oYnLfqkkZl0qTNiNu4pFnmsh9750kaBodyg6yo1TfYWEGZGq+
ZRZ+9I6Bqb2PHrhrp0a6vH6g7z14dyRQ624cCaqCWz4iaH/j7bMpBnKif3OXReSX0XUf98g0DcB9
13B09MjetK+kq8O0HRazT9N0Ko5Edu4vlDLjJh0sqFn459Fdero8RyovRUAqAbwftUdumtwdLG1l
zl2YNJnUiy1B4NgHkltlcFQag5vS9llLfWL2vtWdOZezMC8m1j5rYgZKaRO8l35WCKY9QgPlm4Kl
et15GjiYCfvLOydIP+wwYF0CXJN9Gh1twKzfQKBrSMf2cS+2ylcwsMQ06nOiJlh3lqaQ5gusFD0m
MJMF9M5Jo2HMVVgAitkZPhfPK76/2ayPWRohE2qNpM+Zkx8Q9abr2qyfbZle27iDyhDRk/hk8bBi
tPswd0h+y7GCkY/+eO4esfMfPoGb/Oa7LZlwqwCg2kKPzAG36RhVGMR7UFGkp7SMxkpQNBNyT9xe
g5neAoB/CfgXx2inO/KtguCqc/gWHAchVFdP/c+FHWaNu5HhvvKO5EB3ikDa11cDm6S77IQ0XCFE
wYqwaBr4icA24ybYdqJoTtKlYuY+LZ47nZf8gKceUrEfMFlPhTOJmcbNY9delBtfC16gUshHa/9E
1hqgTF5aqOIpSWk4+GkJRLg9A4KOleQYKKaS6J/BDW0XZmYvItBq7oT/4RHuNgna9DPk5Pj6Ws7/
dmEgpUQWRGAMLz0YxMoVGfxR5vd5/MQ43xgaivmWxCEiwY7BNCPytjmoUXxOUn+AsPXGJBlx+FH1
s7MTpN7Jka5L6VkL3lX7wn84+PPBx5on67ARxptQVfQwt0NAQhQM3aWaPP+d05Kz4ncdRlhIbh8X
N6bcsTE+1EYcs6CYBCYuRJmOnxBB2dcYkR3Xd8/e3d15rBI59a23iu1DFAMjxXfjpehTN9ZmgZ5o
KB5ue24PsGsH21LXcwduNHxuCWomJQiO7EjE+Sqp3R4/SE1XQuoYn2LaPSdFAYLC0Sqk4N6i62L6
Q/29Arvduf5SD0yFcgM4SMWqJJapdSloeJshFg+7vmTeK9acNFLJkeC2/z10p9hb6Jc4BYv1XRZY
LRv/sOL5aEddg++K+1EURrS2yzmSURPnMfMpXsaYKeynLxX6USgnFkTDEE3FUfcSIQdLDZRHVzXM
SxtSDh5rluJelsVdQymN4nOuwu+Qv57q2N7Gzx7RhCUyEDo2jex1gBgK9b9X31dxU8DuUKgci+Ul
tqEor66600R96S9iNlS0+jFuoMgvQ/WmQa2wSuicEZ9FslhKe1R/BUC6xpk7EQDSVNIt9pRAO3c5
lSMsfXIS+T5Ba9p7aoWfj3XLnMOnEpoFF4pstxoRM+2U0KzG4WOsejAsH4N/yqywGKmEmQJ/yRKn
Lfc8rYkr5bFE5VUmw3RzaWRzog3jitZX9qDqhC5i+4zJUyF76iu+8iz6q0u8kNthK4QWSwlnKiL9
YsCMOhw+dT4FQX8e1krgdTzBq9PQTrsrxXDyTYp1zBPJse6RksPG1avXEoTypxV98fOM0lW0uRbv
MMJMvDjke9D0qKkA84TP0ZMfy2nu03f8zrCyyXyCnBTeeLiOGCCJX4f6A2AEBXdmyU4Ried+dy97
rimSYddeA7DlWrS5DC0rBoLKWnULWtGe9+xds0bcSU7tLlO4MA2g5O4JrY6thtyaKlS87oxujTWG
tlxYKOboqpyAwpbFpvA6NeDSi96fLj1MSOwOXjBnichbTer/TWRzwkDQrK/aCzNWMxamheDoPe8a
F4+Vl/bpzfa7nC+je2zTzVSMonxFIaTY3yzjIiyjiDJUmCkPrEDWZWqXyEXp9W33n/U2DR4KQMfm
4TKud2kJUUm6CgkYFxUGAayebrD3sCKT1bdTEkBYO1w1Tk0QySO8HRqUejN5DgcV7W57MxSsrup6
dNsOmR5ndZFJJc9k+sliZSS74e+6I+jfqFvQ6fyhQmfCpoY9IYExQu4RWJ4AJFEr0ap6eh+Di9+z
QDFZ3tfxbYp9ztKRHIoAiAlJT5Sy3du7QMKtPgdo9sax6oyTUCVM3RuCGe7Eq/nm2LK51uw2cbjm
ErVjiUiFax9YmcIweN4RqtPULMRSFwx7y4hG09dIO15aL+Fi9QcudK1VwyproL7TfYn+Mx4vrJce
aVplN0AkiDSGolJ5CNgKs45GtTcP3Fb5cXRBW169Jk0axvnOuZfbwiugJTNNaV0Ghz/Xo8CRQq5c
Fml4guGrD2RVMwBEY9o+FihCE10MBj17c891wsdqTDiMwF1h67z0ql0ySqJZpwtE9VuqvgaY+Ao4
HhEYCJMVh3Ts+OIkpM/KOL73/gyAhuDYgdZPVjA8X9TEvKRsMDHeP+X4hEdM2IPSG0ZWy/TVOxdH
wuPcrnBz0o+HGdwQ/T/qhqCK3wE9ClXElZSIt3FBHdZO+aGwkEW5bm/I/+jo2DzdFi4Wlrm/cmPX
3qh5Jd3rjGdHI4PN/QMLC8OTzjjHReROhRns9ZPCyNGMdiJULiasHzvBoFdRjAN4LXePAgyPHMjN
o0PnxUXlMlE/JRVpp0dr51/wAUUmqntbE7/vHuRbv7G+JKA939vZPKKaCVI8nnGGiMopHiNEjdGe
YLokNnUWV3lfcfuzZ8nAxvMhjSokyk1R+ZgO+cYSP1IEEzpmKEEqoe0ik+zX9a/TGypA4n5hATUj
uyJkBH8f14ixfhGKHCOxd/hwLQRPNELcfYm0eUzGd+I+U4Zo8hh0ac3TXOU+yOarzfslbHu6rmY1
7Z/vlESAoyXCAyyJ+dCeI0M4CKVbIqcHzUKtKc1+LN/QwfC99n7Wg24U526uPCYVDNprUN0M72CL
6v1jD3e2bbjMfMXvqi43n2pnrpA5mT3CLbaJMhDIYSF/7koNaJ7YPRhJsMHGdZ6Lq+wm0Rgm/2Mv
vFgIBVOwKE4RVcr75S60+uvSlU6UzWWRURwJ38xLgNMsydiv/hJIbXuuBmDQDh+IOjFQMHOQWd2Z
zrp/0etGjpdS+iEsvg9uGM+tOIiVv+RpN7O1/oQIJZZh8SLy9V8rPENwIT9XB+0vBDodbcBtT95w
Efb79wjaaoSRQAo2hOqZM0/+GiCYx15xzZV0+zVGnQObZn1KL7mJQ6zQkGYuytN14gVD9OGJu3id
TTykKXKTYzetpfWXCjMFQefdRTWOXl7pfg7snfySBHWX+lH7AVECiGQQGhyCf19jiD3I49c+jU4S
UbU8AXy7LqOuOGuTfo2p4o3xisA2VaEO093oQjNYtSf/SgYxEM1d/6EGbKEQC7RdX3AN3SQ75nmK
m934ZzT2X5f8nisIpvlvnosQh1MMNtTg+TT3jWIiunn/p1DF1eVwLKegvSrkM4hpAq61jDGuiMx2
E0XKcCDPHSoAoKEKSmLdXvGAL9jU2n/dLl6VCWj5OEuOQ8slBPzlASdc0iJJ0zuNtWLA1RK+k9V1
edpo9CGKwdoccuP5YmwveXQH0vYYNhcZ9FkR0qD5WQoisNNRFH+rGPRzw6W+dAtWT/pFppU6pv0j
mgVyxp76BpPVAZmyZwAPoWEKuHDlOKC5M58j3gIVrAx0dLDRzyPqCKdmQ3cVX+vaz01mnTAxFYp1
nKwmzCUHtBt/SJt0Oc5+EFlhbHz0AKXSvlIR2ISg8AAXeQkeMXizaN5fZZqZ9uhAZqnrsm6ESG3C
ARY9cuK2goXb88fdfSD0bCE6g9x4/+nwo/lOaJ3S/H6HtOP2PYCU8JzVQRlWgdFVAzvrWLwAG1Dk
LHp3tZis4NaEgf2O/LZE1uogOJ6rkXAhC94Aoy5l+bze2k6xwOg5+fkGHS7PFfOXaiQswQGMWfNv
MqcZ6g3HjFuSt7b/TMrAgwlmR3iHm2hUYoyfWW2MUI2TBAGmTCiuxKVHRsYwcfKJ5sm4OL8pYHRq
6HMWrpiPuKHqMhCg8YHfzdM3JwZcToX1h4bUGDySjFUEaNmjiIPq/aqCHEm3k1/Hbb2Che3Tw6Rx
TFDHeLBwitqGi4DBYfUNtLJsbfvn2lPqD+AKpBvihdSEWoBiBaHmt2Of0mY+8csj6Ndw7gg3vocG
X5lKLn5iSX6Gau0HiDbeiz30J6mNx9aymhuVjWsu+PXlz89nwAxri1CEG+N6FwpruT0JhIqG23/4
UHlhdQ8GyRBC7Uo8UGMzP/dT7COzr1BesvGoFQ==
`pragma protect end_protected
