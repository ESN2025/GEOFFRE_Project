// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
tHCZ+Rk0tMKuIzmo2OrezYiOzzfLAPXkor+sP4/012UWXsbLXWunvzJNRu4BWZAmKYWWKkTmz6/k
8r5kpWIm9vx5p1HnXjBUm+uttCZJs4FFmDAZpNyjGS+8ZkGsHMJmVUkWeNBQMmkENW8/UOoXQq32
ixKHAWq4ei33C5dKD7zUQuhFtU6lRA6LMb8Vqvv/BTa0t69ASJjDhc1VsvPbCJRlMMSX0b8xJmG4
jGCi/bw+5RvnRl47qM4IHBPDkIAleaEcEfwTSqKafehbzRXj1Q5onnGoWDCTi+i64u8NuD97Elu1
WlvcPwJj//B3+pA11JMZTlXdbuabDLu1MqI/lA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 124688)
zA8XFqjCGmtCKPx9FFLhaEVpBWAoAURvj/Ojyfegg++2Z5KdyVgP68NpflgIVJdBZX8jBCTAJcvD
snLaso/Iw6Y80av+JPY6oHr7HKhHhJJnYaq6AliuMPnseoV7yiXEvYQQ9rQAjtbGZDOsWC6zy7ZT
Zgv/NDTXamvCw1zOYkwJ3LXSSUuOYIlWRbfTsYa5zLR/+U9XaT88ZXewHZPWAlVPEYppDUKj9OqG
z6CcoJtohvBPlOg878ZszdYyCrCbWqoslDf9wHz+3cooSLMMR2MPGMAGQUPhTV7GkTXNg4Va+bfW
4ZdjlIHI4H1vkMUedAHNV+3LVxm5lxyk80Uk2nJdiqv/DbffRhEU1ITAhs6ZFy6bBW1wk/7Cyoin
58iEKudFbT82yVX29IkKZ1oruBlQrV1INZDwRsBAdi0KH2/RLO3X2VfU/uM66mvQOMSxPRU0EJV/
YWLhQ3S9Y8kGqnFHG5M6ZMLGN4JgtUO+Dz7Yev503jTrx5ekll6mpFoHSJZ8j1GdqeEr48Hcv8Ed
XFVo5rRpNLP0L0xonccgR6HZOo1zET/1Fg9Q+BSD6DBvnQ641/m7ccLeVIW/deVfsc5h4yJIIaXC
cZxRBFjqFoMN7PIr1bPKtWNd6ZU5AULzov+VNJuVQpQUkUOn5tWdjiRX8dTQ82gxcA4hMSAiUi5j
TExl+H2LgcOzrvzq4N2agEJrOkLaFzY8aAy3NuJxJt9ICsHgqZM5qh6TABz9yj4J+boBFORJFpHg
Fp9pp+8wBqurb9FAWTLUfOu0v8pIKfJW6tsHF+ZOWQFwTq2Mcqza/cNC2sQsphfU+uMEkAw63NSp
cK6U66msIzVzgVCgUfhOnu3CGMI0gqyZJiphOoFUQQbXCqYPcIUJUjPDt+Hpwf94C3hjsXkXFVuQ
mK3n5M3SuT3Y+nW4JPh4ogIuqw0bSH70fC/TzLVtOqMOHKhe0Co6jUGXAfWhmAFSLASAEcEXayAl
9HsJ8ABne0Jj/7rYBQ5aCX2Cvuaq+mOiI6pISCpdc5xA8PMwLAFwDR2hiXjkW6Jqgmz9P5wZvsLT
8lkVG01JKVDteZsvKgA+5qxfepxScZU7KBacQCK84pA7jl2a7x6kgJLrdf7h4MVIUBaQEHnCNvcR
qaDZe6zni6Ivd5ljjU3aKjsuQ3HZDSh/YZytX4K4PSTBgDyTYClXqa/DPJCJJ/zX5qlOeLZ9jW1Z
rqeKNuqq17es0GajVrgmaBXRBAp06dA/kurm4+lhDfgBTV1Omh7QHtpGGwIzusIaHq3I8NpLXcW6
F9xHPm2E6lAC2joSYb0kSsci4fgOjw2psH+R3GuTlNUbbGEWHsS5uxBuiUvQ/vM8uzDHMjg5h8Q3
A0+nd82ZekntIkVp+ZLB4xqjo31x0ammOfaMDQ2yCTyTa2tv0XFLJNeLyCGUseWsObPWpaYaDV4j
GUvihnlYEpTS2tt1bReBPbpsmggjkRDfmMAggEAauNC9/MuJMuSLeTiWyc7UoJE0lz6bqi0pv63l
O4lVieQOycpJn1091gZK6PWHX8LBu386bJOVKEBXJBxtlesv23tjq1fPdtA9GjsdYMCVu5A7/uNy
sXCqAbbVe7+J1C8xlxWFZeTOBmPRH+tQ4Sf1QonLSsu8nO2a65a2szL3gdbY5TSRts/vjia7qwhs
Q028lxLZSRKsROVlZjZvtI4fxKQO/v9EnV8fxO2MbcvQxdxOHdC+4dyaFjg3OOdAuyaGns1y21FV
5vfwTpq5mpIUMyLrXmci7s3xyvz9kblTI5HKWo6Lh5SDM7Zxgo8iWJS0D6bfuynwBjXDLew11RMM
9HsHHZ8PJcmc7vV4V++iNeyfchsp+p+HQnT9a8EAX53Olhv0ge+bEtvja6DmS2yTgxOF4dz+tRps
avPU/hmfAmu+09CWSe6toGOFO7p+pqjnJikex90rYXxnPHPphvmW2T3WAiTfvZdMnylCjE3l6y3s
CesTJizjk2cd7T4UN5uiCaXgYyXP3dHutjUjV5GXl7gaWEFvl3o0friTzG1XLMI87a58+veCKQMn
3H+gGDe2z40myvHfWO6bfmpUO8eM8vTRvV530fRlzzm0bFTBTYppZU6VcM6jxsJeM8Ulog4BDc+E
IEOEPuEH2+AMFO6vXrdKDFVcvD7HU2jqeBS8/SH2lSo1CHtgOwAVg8Jg+MpW39PiuXohxIKIX2s4
sIizg4kyxRlHwhep1dhN6MG6l3TrAI+AFtF3YKXWNCQ+zm7rQOvPUHKXg9zq8UWQlPNYeAPA00tG
aK7VUBjL9OQYojaY5CbXL7ErbySnAF4dV7qd6UjXk5eVn043bY/jVcU6wrKY/UJkF2+FqpH4XVKy
Hru2H7whDQruksg97tItKy5RU2utrjCHT0BR4NIRJbBNH5WbZGVhIXofK68FqdJq59nQS2q/QXA1
dNXvrk0oRwRIR3/13t8Mlouw76D6oZb4KUwvKhXWl05SSThHiyKai5HiJC77OI5GqmDJD9uwkz5c
+km6OkdDPPoI1RXlKTkB+WHyCmC3icc07wwqVbLqM68VyZRAvFmAJApk/vXhiJAPcbPQCgyGdGHQ
1AVh74uyvxIYvNGI9IYKAy1vcqXe3iqy2lAAAyvKxQ+3Z0DNpyR4O56Ej03gPqBhTg628l/7O6ZY
x/5u9oKwfzwQIHqo8znXyT2mQz/7iV226CJfhSWok7kjbpf9unzxV0HFL5LRMwJV/SY+KqS0GBRM
liE5rf/Jdn15ppuvV/UfC84Y09V3PvvyBY3xE+fjF7R6H1R8wgK7rWb6fppdummqC3EX/2x8jsFr
nJ2mdVo4E2wZCaP1fXOSIL/4FffByu1E1yvIex3lEQ6IOdtFbl97OyNmXb7foLh4UpDh78Ocv8Oa
73kZn41ItR4pgwO8kx4IjpkNT4NSChxBbxaPBmBhOI8MAjPKvM0jOqH1JN6zGwho49jHGJpEg5cq
yLPUL3I7dRRZL7QVku7DwWgtoZXlLsQQiaZwP5t14HKb5DQuUZvhbHJ9+n4Y3ctWPxNqlSLeA0dD
hhwqY5iVHytaTRRaN8/E9Y2WaKun2FXy/GiBJvhM2FmHNPIvZ3Kq6IVkmPzuUhIYQ+D9ZX/Q+KHQ
Atlz8q72hPMiyRAW02VBm15BOTuKrZS4AJTgxHzxHdlzXjaLfyVdOtlE2miaea6xTIQu1KrwjDG6
qIkq55LFGqdRssExuYxTVouUVzT7DQ2rvCTeCTXsZGv1hfwNHUSQFicJJQp9H4YPe0919pvmIbWx
R7JFDUCo1IPlJ1nmpu0TmlGYYXN3amY/6XGEqJv2X/WZNeWfn8m/DdyJtcWxQ2d9yL/+E/uH7I1I
43ffgjS6q4/6GsLzBq4uDay9wJGvEVNY4yS9qvLYZzIVbpYZSUR2X2H3ckNcXJysLrva/eeiVN9j
LLLsz+Lukx45ofFot/maN8ULiFBKOzbwT2gW1qa+iQ7FTXntqe0n7Kjqqw48N8iDlUSRjnOAoZhh
24LwywsGeqW6lQavo9x2zGCLy+pSsf+GzU0b0RFy2lAtzue7fVx7amJNS6TQfI9wZGgMS6L2QUPe
WQY92ZYXlR4VlTcaagCOUMuAdIKwzvl6JFW84XG/6eFOK/6+iG7FZrX3dDj4NvMYKYC/ykTnGin/
MYYWm3YAP7SuVnZj+X5HFVkBc8RNZcNku5lb4m4W2s0kbIGqJptr98nKIz8eLujvV5sIshY+Mj6E
QMMjNhqEEsVa/KVjkm4+WrfiXHNH/wNVMnzOc0bMjP9TC5DXI5Ayj9Vlp6cZppQaq3x7HEpyip6S
4N/uzrvYYViF7e/ydiRgGagCixKdOjwrW2WLzStVM6/d4mDUGbjJoa3/L3Kka3hgt/fnZiL739ED
VX6QtRWmuRSW0Vvl+Fj4zc8cHUG/0xInb1qygfUTOXF/YqzeL5p2567EKuR7e6UrMYhsuDkDwKEG
q5kuRzAnB7Kil5wWsnQTYEDFlZM9m6BCrdxtjFIenCzgLojsIXRQnLkuJf8cWtD1t6u1ufcyJe6i
cBGJDz0+QmEhBlRucG1WRxf863CpadEeENEZTDlorQYZM+u/cDbKK0CmvsNOUhPaVE12xuYxnKWl
Jg6y6KBddiQTJMwj6ZZhp6oZaoWqELGLyrAzkGThyYIDuLQc+bywfus/mtbv47e8cPH2y0PME6Su
xPeSNlXW1tdhAkVhuHoWd2Mi84iMcGWWeCdVTwGQJpf9bbcjlL/dliznTxqwNRfaAr6tw1u1Ki77
uDVRnr6sDj2ookXQqwE0ttM1OAK7Dt6ER7d6lgLnCW7NoOcZcnvnaSCYt1/H2neYxbz4rdPI3kRu
0fYwDlZgOk91u2+N+XbyGUWCDrG6CUXlUTLxR12DWflZtQBOc53ZSXyr3aTcPqXON1upEC1eD8tc
2/lIrFcWJkICa3Q8rBmFWRYiZJX41l76lBcJF8Gmbg4z+9FKVmDvULstN1YZr2y2PRwHPqyrDxUD
Kp0Cc2FSI3sMKODaAq2Xz0MBdUuaTeGJtYxSdjOl+iP/OsOdSAnLN3HOrKXAR0n8pz3D4nsoVMFM
TRNDhBxA2qk64k9c+0D/9wSGIGylJ5AhNaPiIZWabPzBROJv47BXdy5/T6hsRhH5YJpD9UouXjiD
Ou/O90wz1dDYmQMT9wpcY/O5Nr0dzIbJ6P49elB8cXzcvoCZtudEvnGMmCPOED0JOwUwMdIEPAwT
KzwOQ9GRZcAuL7nDh4w3Rd6lktqlt9R5M92cIm51CBpfYoth4vZ3b72S3vjYNXEKWSHKnesCO0p/
WHhpQyrKHTIlvlFJZavN1kjsH6qd3TS77O1Z0+YoAVghAw1t7OSAncHykvP4UAT+x6PUkz8i1s5f
Y45Doj6x9xlLl2jjSodTA5Q3o7JuoMpJSTxMsLx2tMRFvbslaOdIuAiSjeOrUyJGJwbUeCBEScQS
tJVlkJLu9m/wxm2m956hNIyLemuz+67TvbJPPoePromApMBivSRhSpzElGV4FPfzufC+Vr1BdS++
+f9jfAsE9W2sRyvDKMSGRQk8ZahosZ2pxXwyMtuEjC4UONP+rWFOXp/4HOT1WYldyNrfp/znKIoJ
5HsgN2fznu0LIfPPa6jcukc+vwQnnV8mhqDVf+cWe5dRmFTXODjr4/IoE+Cov5QoroBniDZbJ8uj
v0s15RxkVLxKsh9ebFPnKh4rR8WkaJtUlsm/aBxyOByiRj/7495mSVCauto6SHcRT6ijE3e0xOPA
+2rKZrVWKAMCNZLEZHZOPHa6n4GCH9La++rj9DrMY//RRJ5F7AIQt23z3Ijt5waKmf5IMfMfLOKV
hGa/asyFKnmaDgxV6qyKvOFscC3iYOfV+B7MUNyeAaAzzVvNpUIdpssbHd+/LBsOzyUVtN84mCIC
HeHomECgRM1/2MZtsE1+xXQ6X5kmHluGeUyXPEpFKY1wmMiDsXOozH0RSUjb/GgoXwOYYrDn6CcB
wAHJ41uAU1UJjboC7ZEiXxbxa6brdn1nbk5da66G9t1nVtkqtEB206jR/axbQPtYkZUYkyAPj7VU
fB+xyyl0djKEB+2FIUs4W9WtJBIkqBHIUm1k3XQo1vK/UwfZhHVdLX5E2Bvq5ueBoVvHrH5xwUvH
C6PCUISyF6GcEk662NkiNaKBBI+hADhFUG5hxGqMqIcBl5uPfruM35tsFyWK6FhaoWiJuccAIhzu
pkjNtjtB69z93/qsQ7Omg91RN4nVjHSQa/jJE71xclol1csZ5Z0+vK19hciyyFKOGn7qOv241MF7
3f6X8Sotz6rpGVs0wBi6YsZwSifYRqvy3qR5w0OrmU9jCaXHT55HaLbcANALRwm9svVxPKjqj2FJ
N+fvpuAtp+CKjopJqUtcqFjEArKPn3qsWnJwKKvxq8f5D+nL0zab2C4M1P/vjLnd0et3AAYBjkw3
hRvZBXh8sK2H7Hbbu+XgALdaljAPnxDEJFgaOGNlk5UUOVoGM1R/MljH44L9K4f9BhrYET2Cesqj
15qpcycNzVE+YmJffzHzgABarjjDRbfEnxUbTm3uNmUTXhx70MiMpg5gJ5wJwkg6YeCZZRzyYLOj
bwbkd9ekabcjrT2C19+4JQJsvs8K6UA1s78GuMK5Jgfzjxid141OHFzSF5Q3V4NGBiQGRXU9rDbm
roXPQG2afhRF7ILd6Q8ss/BzThUXRbNcUQzX7N7/N0IbT7cgLmR/E5Lt45YxQJH+7G4wpHpQ8IRq
KJ+ySGc38aLkBW6cQk3bQ2180lhjb4UxXEWE96KaI5UWCqAJ1pNCWlP2D6ej7etjYug1lcVfkl6L
FmJNv94h6Hd1izcT4B4CzutFvHM+RI8MHC5Ma1OBiAeYBS3ZwjReZdKCR+1ynRX9CedkabNYbgrP
wo0jxdTRw3HY/2KoHWFMO/frVaxsbJmVgNBvgbzT7dmQ4My9V4v7UEDX9+LDlO8wts6nzG5Z3dC/
L+HC7n1Zn9R+IjkETLtiv67D0mY5xOnmn+3IYslmXPYQ6R9qqUGVcoAcItd6XODrsaOt3k7j9ajs
cWDpxCY5+eKLgYBkxCw+gDDkxW/45wC+wb11qMkPwJBmRasISWMF74pdcj0QWjbuNuiHq4kjgslt
CdyCr8CgjzsqWZ17+2Lk96pHsRJpaMYA3zvwBnPQ2le+4oxNfUZ6lt+Zn0VCNJd4H12bYzazSf11
w+dNoYXKkSFX1Gklj2BcJ0Gv5MYqmKlEsHDNzz4isI7eqJ5O3Y1lg0diAJj6+cOy7lWadde8/mMr
eI4jPrtfZ/mTRvNv7c58Xc4zWNZW5wwvSuNTlhssoyEPH/11ceLPLwAKM0S2emiMRUCBZAioLyTj
J3IkaRPNQdV7gwyZcixaVf8oDvxeEHU48uN3n/doet1ALu4H0N2oRwBuGOlMwccgE+IGETdKu4Ep
ukUl4JBPGCB2fbei9BJV1nbr6jL3N24yQ4F61FDU6iApCBZi3BNPEotKyqpzkELDPfGkPk9CY5pI
/+z8IfGrd2EnCFcVjRjf8/esoBRtq5o9VkJabLF0NpTBUcwYpjfDribfGxYMuOQnc848cRyEkVdy
SMS9LY+mDsoEuwGosNx/n/9Uoj32LqMkXwPgLooYRP8nWwd5XBM0IO+XCY2wauAxXlaSqIld8cHp
+AKDDrasxbeJd0x8p+DIOXmsp7kW29LX+tMJcQLy5JurC6iJr31qNUBKaJ29YwjGPec10YcMKpvI
53kRjUrDpSQla9RoeZ9i4D0HpQoLpz9+V5lOoKNLpHbSF1UUWBmLkELE9Nm8nUgGJ8MXj7Oy2+Km
lR2gnTex+GOGQFEghJE/MscYh72NvvDKI4BnAuGH/nXeOwNJhz2/DSALL3A5PJYjJFXYekBs38Kb
oX9ll2HA8iIsLT+/k+TfRLIpwPcFZ8mNtqUDioUOV9TSn5CIDJoTiBh2bZCCOPb83CfYq/O4ZV6T
D5a7duukgcM3bDyDeOpmSwRgPjW5Lg34EaxGK1T1RFSygBOF9ReFPp8/IknX6JfzaXVVj6dnTnz1
dWxiKzDIcKRF21onzphNPwDvQgz7rtFjSZKC+pujWdqLzfkJ5AKTIAkkUkwpvZMgHUneZtQ9HUBN
okFr9799iGwCFbZ2krdB/9QoTfoBakIAJ6QHvWgEK6+UCVcHdYZY1LAqtSCvvOiNKUFJN7m0kXRv
HaM8sfuoCUAXmp3y8viFvSa8RmcCkgBmjaBOVg4CUF10kYdBR15SemmIiP6twOj+7meObfC5QKco
62ZedXa5tqxQa1XTIMNtdfmzbfQsAc+Jwyv/0gR9v0BpSfLCUcTyeVmiKmpWhRn9SC2a8x2D+/vC
UkQqmKpm7xCPqUso7di+HkzSElVUrl7+PWZD26U4wZprmkwm97AdPLuayBIHXCf8r//h6OT0uToI
+f6YzrLXf6qCWCg1o2R+b8jcGQrjo3yifj4LujdRWTPjeTVSpOSI9q/WzYDDN46KB06Yqsx6k854
I1GWc4vXYdpAA2E6p/EBj+sf9suAHm9R3EiWyKN1paz/uLGyawmzcWJ95u/bU+8VBSrYo305rUAF
vvT9isZ28JinAY7pKH7ercs+I9FwP0zpYicOBpj5B/o61CtoFJpCyCrFZqux0cpzw0bd8UeE70Gb
wpwNFGSsdeMfvfcW+4B7ExcCEXyXDxJn5zjI1FWr+XUxg0PyGYYkl5okDraJCGL06nQ1WCk+8kBk
W8qA9OMfSR7q5G0WhqSffFz6is1Chmv2IJhIteNmDbtBQGPaLSQGwCXkDf3zS1K9/A8K/pjyDZiC
VUxI+DwLcSo9uRQKefuEfC2OIEZT9OP9pZai9eekIAvEKD1I57jzqFmDP9LoUlEVHTAAhVlUqEk7
rikGCyqCDAMNQdDwyfnE+snO4DIx9J2Zlm4t2KXuFAL6P2mDGJXw6GqpyLawo1HX8C6xpgRctqLE
U4E4rKgiXg2cgpnYWHmSjgVK7F6WI1d1F0cs8CVV9+DhcDpwSKU+7PKbYuBkosRnBZjuLHhyt0Fw
TDsDmRku9k/fO6hmcK6KnuWWrSMSVKBwkJwLfQgdYyB6qCWTjxO8dZIldopdJF3P/leCeQ7B1Whi
uu2gRYcjJV4rVG1VImnj3cLGI2B9J7jlBOxuMxVFX1mdxixJjFNBTDqafxLe5iKMpJ7cIcli4vkw
uk3YRd+U2ybPjtgP+VZJQe++yPa4qmG2+L/PW0dWD6ROcQKi3LVGkKglFhL4U6+16hDoGesqmTG3
Pn6PDIZRSoUTa/WZysyRXpVgDsBTA9XIob6m/aWkFkxzhmdTzMoGfQ76HaNeIQx6q9XnlZTQXWpC
ZSrB1G/BvQdoU3P+fl4D1msSpy0IM7ncdZw90cnP7w/X5ZUTc/1R5ZSj+GkRGw9woaXYPtYzr00v
Q9Q4TOnRIAKzbAUd8Q6tBPzeZfwtLiBg/5SGqfWUM+hlURoRdX9TvJVL/Y2zF2SybAin5fx/DQmm
nIqRYzNoywG68QG8tAEO8WlI0Q2JfuXXfb45mA1UT0F/PoXeRFKgI8UX7aS9sDGLisElLx4fiu4O
O7Yqi01jlXW7N/QEPSdf3aYfhAfZFiYJvgjiuQSot1uiXnwMnNY7DU9R+lCLARj4wVZXoYzBGMv4
icLYL033qrac9EsWFXSeM6qNfiwZXceVe4XYkHmDrj0396QUm5Fjto2FELEK972oya9wMUU3FgQp
aqEIO3kVPDVCV+aTcOgcxP3OsQU4oj5IGV7UwkCVa0Nqw8Rka0u38Ky9+XcQIB46XrQCuBdknXpW
KUQDSQF+32Cmpc67HrTrEhpbRF3Et37C+d0Raj7U/1XW2cNGmNYbDfVOxr+Uh5BvbAEKBIBR2XP4
ptocvcJX+jUBYx/nCh3vRfWqBsorDRfAMtWUHtdWaVtcGX9jWV+9adXpVDrVlVbXO5VIx44788He
IJTQ+K5chpJmEX0JRS78uu5IjqcStpLGHRIpasM5KeuQrCoKmjoezvsNJm6R58kGj2HgRUjCzEdE
pMmxRb3rAflg5pMFK/hYolDPNiY+69XiuBxwZuo1I4aQCQLOBGO3/7Y5R8heZ/wr8PYw3WpIKqyl
JKABAovCIBrYBo5x0gvusqIdNz2ylDFsc6XLURfnBt5csN2EOSdIrFuY2WZwObpNsIsmidFp63cA
ZsN3TbHfop7EwFLcKTrhkKzudymdAdQmHs1B6MrHV4BPUcbzgnbyfIEdodUNIrVILvDcx4L+J3ES
Kw7CxPaVSFe4edYKvFv1IKYp9t3m+TIOl+6NZ+tmX+0aTn03yLAtEyKmUuLCZOyTYx43oATFWRzE
m4YCGYZ1ofZUMMDkNRjGVlHDZmodeUIbXVghs0tsJLAqmtSmHaVcf8iFnzDaqIQaGEGRWGUYdiVS
8aKXrTRCSl+RUkMoXssAX23AAatxP0WA8muuzruI56DJ4QHIvkqDnUrU+SiXr6cqCdgn0fjiUPE1
h04ecEkUd5zoVyiBfQnNoojrRf4eRmpRTMVYF3T823i2W9QWab7MiJKfAlyY6tstP0EriGMwiZM/
rhtP77JpFcsw/ou9PVFjkpD/QBkl0apnZGiGputtw95mYpuQubrQiOfaCGtuMDObU8UXlX6b1BZ2
46cZUs1O8pvc7SbQ2qKane8Zmgff4nZXPkfHgJfxnTDaFS5AXGwg2rKNVpZ0XFOGe+t4RNLxXd8v
Ex7dbVc0k9UPEP+XXV+nZrS6r21KHVza5r5r+LIaW7R6fXIde4JMY/7m+Waa1xLn9aRkJC1AB0ek
YbKtrdjk0g8/+wCwc6sqMXlTI51n2RaS2EdS9O8IwrGi+r/4ZWCBf86ebwcUUj35EbSDpotqx8xI
BVPUha7EApY5u92FvMwUJWe0/eTSFt3ZXQTrdtIQcKm0oUzlhTthvpG2+OLF3xCxf6hO2sFnFouh
SxmX+9OEz60VFJLjYWAsCuL6Lw9uiJxfNMOk0zY4el/50CaLAbgfocT6NyqzxSEq4PfNo1c4akej
lv/2hldaJBeOot2wS43NC4UlwBasEK48DyW40ywz8M8NzjutGO/OWJMaKMxwMpXU7MFA7oR/5yAv
/V68/tkx6W32WeKEQI2lwWPljd6lobr17vrczV71iCR/cFGrKeSaO3dQvYW9VB/Z8Q93SWeHINkn
ur3da7/Q7CTmHWodGfMzHATj98FdIbrrjUUv4/PZd4NsAsKDauz88NgGSRvaSDqqMU/tCwG/ker2
1rI4LqzpuPxNfIDczhdEN0V9i/Wu255hLTWrmJMCEtw0rt/7HpcPJL4gkW2WkhWlS/1HSuUKDSdZ
LgKOA8vLWAdBEJfWLX2iiJ2VPD3fXm397ie5ZHJ7Gmr0IzbcOcveX2szlqWPa2a64FitEjt3ACFS
azU3/rEIlU12FX0McGk9yPmAAPrIN8IWIWmigQT8SCB8W4c3Wqz6Ri9hOAdz78AHst4GQbFpYz7o
5o7HbFEqfxTI+UJ0Y1wC4MBJLwyjSQRdq7NyGy7a+VcRQY4vK3zwPn182b19/K7EGntai8WuD/xS
1rIcUA+RSo1P1bhJLDUouUtjsHnvIw5J44ZM8UvFXIlRcte6/HxuvfGOZVz9x5xGwFD+KBHPnlv9
TEDsoYfOp5FK+p9H6T9hJs+pRpDsD82+G/nLd9JGC9gvlqGL7NHvpYb29CJf2ncOQJXjq0afdECj
T/28KidlNJJMm3j7IZxB2rDT9odtwhya1qF08jCq3yii2YWOhcA2FYC2YohypxozYy+3PWQHCfWX
lwjU2fOs1Eiz+QwHe7dN5Qxn581YsADHiPvfO1b4Ecxkuoxg6yGclF2e8VKWwl+vkQq5EH0I3LQj
Czqgof9po39qONP5JBvSFQb4/HpIlXNSFTxpz/QBc0SLL1FQp6s4omZw09/odjam49guyUTl3af5
JHDjP0aTWX0qvb8dwnUqDQeVuI13lBWQrS1zW0NcGmH5stloYAra/1vHlmZRuUbw0AEgEYG/6q28
lRRTmBeEKkGTMVqE81meOqW051tDAix1xEj9lDeL+/6aHZSuQO5MD/schqJYGV9BaTX0xvbWh0DO
kQz3SFvfksenRabL5I18zG9yhqclHwfEVWcPudI4UcZxfP7HDvgyN/OEtsN098X8qmohxMfWGh4w
AeZu610mW3/vI0jGx7t1y5bsjaKZNAmQlunZFZoaDY++nWx0+JiHZgahhUXVtXotZi+A2hTXexlW
2sZtESLNnxnmABdStzIFzdDLDWIOERFvY3PsE4wU7VaMEJ6CoOhykWGc5hiyvlSE2H7S+f3hU7dU
fXYHRF5S2E1Hdg4y2bVbwQf3csHV+kaVWhQUAUfEb30iB/WwNAM0fxpMxR8xik54Qvxq/28NETP1
Xw8wqTS1sOPObGnBOPlucqayPE8dD2CQo07zDWkuJiyoMoP2gp+lEAKRTJrZKTuNG02rWW9LNHdi
vxCO+lvVckh/yKhPt8cAv/QCR0ePeNAkl+vmx0h3OUckfuJXzOIl149Ca2G8Fkcblllb7IR9Xs49
wsBYbWVZbX4U4+CulS4IyFy2jFy/NTgJ9oOfjHqbnp8oP4Mma6iCHkJm6kQlkhzO62gOc/XQ1M70
xwCToqvR3RPtFkvnYLzZw8NLEbkbzMTTdGAbyFTBYIvfoxOJbdrFMJnlnqA5ORdHZ9cipadthmeI
YRVkBlCDefc/F6+UhDoQezNlrNUAFZd9UtHj4QCPmnhEt6dfhNU2K+4IchPI/0Kn4D1xoMc277M2
KGlvg1actoVVHVI+H0Dc0KO+k/UpqYYDcaKipH8t0uDLzKQN0vE8+7gL+rHW3FvpJ1hlGvzVc/E4
wDObOFyfzUrTyJ2SP6oInrjSFnLVa9Fr32adHcRbyjAkjN7mjl3udwY+gr+FfIlJb10TBAEDXVCS
T1ASPXnDGGCcIZt241zdtD+U+93hCC/2Zs2p/eihwJ5AuLXl6f6kIDnFTLb1KYe9edG6gUGqibAr
O2Gk89Wm1kjYnXbez5PCrH1YrkXTry56fXlN3Y9NgN0PosKomZlb5MS1S/BtQlCS1UA4R9z5Fogs
uIZLlRWLr5qTM9ToaEogsn9AuNvcgmdGyAeJNHnSTFDloN7/Ntf35/WWdJ//2q2mCj9jRUjMy0C0
weAfE9KiTA7XQIxwGj4V9gv+h0yfxqyA+oEFCM+GiicVi/4Xf0zFPQXg4xQ6Wrs3XB4h1ulMnnDx
hSf3pFNLNgYXnlfkK+0XY1LkqJXc2W+lj6zaA0X0Yq+frACKqKySPiNe/sHvYJK0merG3iLg+cNx
BXGMkXmLEM6JuXV17sqf1NqmlULtdl/lGtWWzaAOU6dFjZS0brnXCkMkMp6ZOVh0RXVL8Jnu1cg+
ysmIDXKuoAj8fVzGxoUj8gpP6o0q5epc6dmnoZSZ7o0S5bKW/b70kx77N9vjjtDvFvNV58Uuullu
xEpktruz/qxx+E5hHxPXvMlWtukE9DptJi98JPA8Ti+Uav96Mdl2FC4VfBFpBUlTLhYXEUC6u30X
8YLw1RuFU0xd+EidTcKvvx75Gr7cm0xON7gsZumQ76eD1Wje1K7wYip+zcQY24Lu+L/sckMf7jkL
jYyt0mS0NXTd0XaxVukFbLtOGyXD4tWU3xMXnunB5cTFvnujlWg6oxbSfqWqyTRGzvZfc12gJ1y9
xrLAktPW+cpDeHWgmd8oIBcgra6LNAjblIg95KjMAG7tBAqMVlb/aCMWZeEGT5TC9YjRYeW5WTh+
ZFptvFQPNHNWukOFVbt9d/ZgNDI8JTXrE7YcmD4ld9dtzpqKnbdHySOIAahqSGBee43Wigrdpuw6
xacOWLZyCpGwb/oPIAMVPBw1a2f0wobebuH+awW2ZgKbSiqPKY3HCQzEDWX27rtrxF+C1GZIhZNt
viZJAQPeydoVmRLdgEkK9JzBV8nvr1nXpCpSDt2RuCducbwv7zp3cUd+N43s8wiaqORfXfdB/siR
Dd2qK+CvficuhywtnWQRjcdWYdj2QWeAUiBW7mAld5Fi8UjlRHz0BT4LorlN+c/O57mwKCq86IP6
2DkuTz15IQ8jR4PqC7wqIK1QG2B6ejspmpVSkmgItrTLo1CHxcT55Lrc6YzZh10cOv6Aaq0C8vF+
zKSidW0QHoBhG9kZIuVWyse4prhTZqOd9JDWEYMEt+adzAShs+mA8J+O+J69CKTMc45ryHrQSKxg
mSme6uyr91tjgtblVA55cuieHCxnlFQOdA4bOAzF4uES+yyEZ+DF3r6KghtcP0NG3Sh9flPbmr5L
UdciSfdk0bv6QP/1ACEi+//eb0g+WG+W/TIAldRWzAtsIykaUgrUTUQHZVt2IPfww1BjeINwZJTn
WD8geYHE6XIuU0NIo8I4KHLB0m+nhFMm3stvLUyCPmFsxXCmfD+/UNncetWc7uRQM1mAfg8VIKA6
NoTyCMod+lK+fbLaQ/GzNvnXZPu/Fe7HvbBc26sSj4rS/sCU6Pe7GlQs9wOYPBYO8hTFJciLi66E
+G2s/xgq8Db2deio4AGKIgZ6R7+msbIqWP8v+pK9qLEyFe8hYYdTo6dUYOEYQfCIc9SjHIg9egzJ
YRsUp7jJz0/dAa+Zu+w7B2mFNpc8H/wUapoYcUybPGzLg1hzccpMj7zBhCI07Eag1+iajzWkPlAw
dWHLlfsSSXgIgH3yk1q8oCsXNljIDJkjgZxvYDM5PUbVDZrWg+/b3X80Quwi6TRXjN9EqnnBZ/KA
bDd0T+d8/rRk5pus0QsoUC5IfHTSRRBujuDoneqcqp4YYDjFbNKjOu/7N7WJsxsOnJGeJ//Rxo2b
zAsYFjEt0macMKb569+YhzNpi+bCvTl48YZvbyg1kEUFukK3LEs2gGUaH3XKA8eLHNdZPBJ9zgPu
8lcsB+H0WmRE1v/ktoeaSab/IgRdfO0f5/QEJCvjL1UhWJKoWyOogcBE7/s9mVLGndfIIH22xy8C
xN7bHOAHaX09GWCxZ7GHPH2qXwFv2Fgx01sDD0E9o35qinI0W90MQOwz4447Jhy94TBYbX1xQ0lv
SLRmNuKtIYLfqbQGSI97jGvsso38edCBpY9Anz6zMHTGW7HbSThl08v/dBSzH/cGR3UvyAZATmFt
ow7ALCm7lX4JuIzDJouBxCmrjYzQqkmP6ot6essiXyFBGGLqRRXhdE928J/GAI5Be5FxvEdCl95+
J3QvPj7QqBZc8D0u5RotFJVR3GFbCmLI+8PPkXCTp69reMl1YAKOe+YuT4WEuONUj7xuQNW2j1RF
5tnZSCvOBEssKPJeKXl7oSyTy0XXj/kdCtFRxdpVSltbZLpB+VQxGggLZbOLbXfQI0ppSKUFIg1Z
4dkkjtZOsqqGI4cwTj23W2AoAiuENfFvMOWdlGRBMm/cv4ollQdfu2FruwhS2tUQVug5ViXi3iBI
66o/fYVhvhmjAI1ycAyY4Zk/5ObKPqV5IA7LNiJY3E4K+GCCbXhmrKbr/vGbvuLag0xK6yxh7FAM
bd0psdnOH2hKsswivzYWseJX2+cv+GhhOmzzJZudNZLKZeVCvw6YYHNts+FVnQuNZtYVzFhlVdEz
fiiB37FfPSPIQwqE1q2aA/cL89xztmOt4h44fTkRieyafj++eiaAMiKrR/xUWwrQIHbYhXv+HeEQ
PxJzyrDF3uJo+nwTyagpa2o404tU+7phHFQW8cAwVNCevI0X0Fyggbf1RkJkFb9wVcwERfwpuPP9
rH8fDh1S9i5a0tT4IgsliV+k9CCHtLSbZivxEQu/BzaVV64R9vVHWY7ARud/4IS6MWjiQJpA/Cvo
x0/vIvbSWXLSDvPQg9hf62ChFX2KHp0izDo18V3EOasxu4CKJgOEKGd4GJQ2tm1ZP62UZ9OY8ynw
2imjk5AEE/jCirvyP0PT8C4d0hTBSO7xzsVXAa4RnQdEbwV72SA4mVq4SUk+v+VfluITYUGspiVs
D95i8f0Kxd7DJrIBD8hRArua3O/o7pwOHMfJ93hv7NkY6HoXIvyKPEIFbODPAERurM0uwwUUqRjw
apqVP/cYPwz6jBb4ZmSb8lRXqBSB0aQNrUI+SBm6vqc+tQIoFLrONjy20aa0/XBl2YNgmxpL4w5C
4IxuiwUyHUPVETeaAhi/OVX/SuQkfoDi9yHXt/6Spbk230Yo0IkOoLdIAescQS0vjE6hVFfW9Seu
0pTKXPFxL6+gjgEcEE5B7vfWZ9Y9DH1s9FaIeuwHjKTR47B59bfkaQlyus8wqWrtZgaNYZuunj8C
CXRzgZbad3H//VR75ZYHhZnfu+vQu3mBdq+pWXbFQqsYiaZYNjTSayj4JXGhL2/6NlNkJKlktsb1
6aGP3THCmDu2XgChIus0YPLEdC/h9o/PhT+xyK8XpINIJoT80mLV01Ue5TlxzN38qYA/gFeAWmxo
ke5Od8FbO6l+eqjb6uNVvR96giJ++LMm+kiQYehlWpX9i5wqXfBsm+DgxiWD9uLBR8luWkQuo6pm
llA0wQpqcAFl4U5RaDg1mDD6lpxh1plfTv0crC7v9wVeBjq2mx6Uej8CzwRXkW3XtqAco9JAqxPC
EbgGkWGTHIOANQbVlgz3UZ3kVqPIEH+BpF2L0Gr9hn0iG4TCT7UmvXe1+WH83b3EpXr36k4YPUU3
yqrme7/Zwxzw15JkGTqUuID63l5YVderH8va6ZVEQ9Cu/9lFxxk5YObTV4WI7IiPQupuHni7FCV3
QfW9MRVMnRVzg806R19vip+CjQZ63UGzplgD92GSAEF0BJHaWTog+RBLk5aRSWYjVivWmVnHZn8X
/dNtuzOe47Wct/IF+IbQ39LFUd5+SHimw6kYhNoBRXNvGl3GN2wuEh/HtpSNCEGUL8cNU2RtKC4K
ndfo540n3AIVcSyoRSBCNl4um64ZJ5mlxP7TXJ70uIMzheo0AiUM6Umy4HFaVhsL9PTyWn/6boIm
OJzAM5tmVmrrj9kNixjNLX9iGFE4Bj2DZfbPv1Kg+PmMp2KdXwNxTVaPqQJLhRaPTjQqrcVCyH+V
OE/aqUS4rhjApJ1XacdiufVaIht/7ZE4C+ZCPPVVxnoRtR1kpnXFs4g4A9XSCxOJ0R6+hyFo8IN2
VmxqddHPwJTgrLlxXERJwF93FzP/48hhb5mOb8exZRidT0ZJLlWbB8lxOe6I+yAHnRoWeDy8yXjL
RsClJmHvrg77QAATOmdCC/QbGqwnm+zKd2YnGAE0M0EMN4quywtiXqx/iBriWWLuJkbnQdHNuxtd
WG6qDePUcl4vJ3tHd5+w37dEqDvqvmJZDkKuAZ7uc6vo0YzMZ3UZHARnETwDZaEa2m9uM05Ys7Wg
OkN8TkG54pKGG7ot4QnEqBQh+QF81Ut+4gE6bvjX6b75fL6XeqhxBomOtxDleQyaR2CQB8eaMtp0
hHEk30mW5GTN+nswIqxfqJNAm8o7bSf+OPxGzGseOFNpqLIAch9+4DQpTavRwPazRAorFX7H8eLV
PwJSDq0+x4Ld8gHfS1KvmfIR902tXRR6n4pPm2zOB4Jp6TOOJSFkHb9tcfAsq4DkqCevFeFMDvYl
kOAI1TXeYo7aIE3+1P5sVP8iBpTgWzT4i5sr0bwStSPc/mozxkfEjC3G164SmkWtBFcJOCpmD9aS
0LKOJdnihkH3148AKE2ebQEjgruyLw4t6aei+Lfj5/7BiGHqoiYRt4TFreIyzz7002eRFdJ/JeRl
JgDw9y/7z/LHm+DhttKwx6mSXf0bTvZPFgPHgNQZWj7GrjBVgtGeaT1qc1X3AJ9aOJRxA051wDys
4yvABr/+qS2GYdZWB7KgWSXTiN4rIoItodqPW/yqevnN2KiJnXP2Zs2rM6r0KRmy50qS8dAO047U
OjXXAPVY+482bhfhutUZI5LRjzbUyIbDJ6poz0DFYxjDV1zMiXhPRPTbbT1M7oA4GgfskHo3/Dy+
zOTxUmvo5kkf+i56yvapMd+PmeFjPDz+74sN6O28FFgJrToUvCgxvqKRl7QhHI0o/pZnUDhmjYUt
cCHk6IDAIaMeQdW7L9mE0+Mpw4EhFOwoYbC0OeANpfWAmNcE7Sztus/zBtRyA5bt3D19+xPZujRQ
EEuQqRfZfvivMmvi5BZ4wx1QICm1SzFxoMCkKS/ukBfJi/PDqDI+CokRKOE7GLch/ayFmlT/kUu+
z96hx4OToD1yXqkco2hajXDxA2C/bUTki6tPUUrXYwa8nbkW9YqI9eODxzwsIU8pYjvHOKDHNcxZ
mYS4gj/kdu6Rfh4U/H4BZNlfvsRcFdG+cNwaVsPkfUe/qiOU2iyv7lzOB2Q6ZbTD/esMD13DW2+M
+Ogvvt3gUafKOLKVDIB+8wtEgSsG5akM7dSo2PPE/CyMCDS+G8o/dKLzwZSlU63eiVbj8AlK72YD
CJaiGT49HcAX7PBmWB3tuN8e/xQ/0BU+niDqvH3uztBfoNgEvduYiLedpWw3bZMci19R2EL7FT4F
/Rc0oGs9XJH1KrSLfrbljlsW7Lg9oZy5hCmg5ck1gZBraNKJnCxVctd3kbzzd7tGW2zuLflx3asl
tEa8xZcaAqljWKMgoKY6qW/dU7qWaiboJYCn8tehQ5ANzlrZ6me1bNjXFihjRxASEuOLjalFgjUL
sUiyeR+AdfT+1NaFZPE3A42QYut4GIogN4M41qK1TFKM9zt1xQjiYUqf0Y2Qk5EasmDZb23M2OXn
c+m5LIXTpx+Ths3ymD/YfWCrbc2hSdz/J+WUj7GHpRVgQvKLm5cCVxRjmY6M4hph4xxk9amWPvH5
RnOJQ0JOgeziLfBWfAdbG7rs+9MlYbWBAuZo7r/DRSRQmJVLGHeNWE3q2RhchBkTYe8D6tAGHowa
zM0y+sDtFOJau4hTOAfSMfjMwQdqxlfc/d+mb1UlP0JRJrJ4AG9YjYdGL/7VYBgLpxsbKebqUL/K
GiwIuw++/eIEiK1U9qAJv4nsEdVmhiI2iKKCkUOyfiCfc4yBK7dH8fNOUTcbfHiSPiQ2kVIZGii1
TYdZuJpZ+qVr0ZnV8c0jhCaSalAovRfENosvBDV839s8LIjf3eIX7Ti8K5UNp0LwC4CbT6xJAV9L
CNEGp6AeKvoPb/i6O17lTpLWsmJ+Wk15khO2aYx0/ghNhFvE3/nMz/MdbiVq7KhSiRHm48peYnO9
H3ENJOQtlvkIyGEFKhn0wSGX6Sz3Sx9DZiuzfDXMl//KX74s3OQbf3ZEtfjA7HLgKf97PQc1TDhG
c0J7zQMh/nvzdLohPdoiD929YNBmeuNwN6JRqFeIvGqnFuLL4kVXD+trHvbmyhmhsT6tgzszgBM8
P9nRtIkjX72QQG0mh1tCtk5x+oUKtwbQG0SCOXs/CcK0GuXe1QZ+dHFZGku9kFWN1hr/NyxXsLt0
aqAqf2Kt8eo6GK0hdeZCiUs766eiR9bKp/smLhIOrhkp1pXpeo+Whkx5EEnjHdoxdNU2jjrxoIQv
KQ73FGKzCuDqeC6SiCGGXdCC0gEP4BRztAHV2yYN3XIN5Qq14hhQdwtjq8rl7vVF2QWQCqDaMylh
fY2DgRRmnwUvwTKzheYxzJCVeMlxhe9FkZzXrs7Djpk+gh9Blv31oq7r2BH0e8yCcb+Z4Wsryx9L
F/n57wnY+zswpVK1VwAU6enTiQhkmRSi07/INJCsIOeFU7InmDdfua7oTYYmSORPd11YGRKUpVFD
kYzwq5wzlZJfuopz6XfETP8LXWZ2zfZF9fqv8iujhMSGj5++ABaw+LGw/kJmJMfp2eeQEhclfLDn
DXfpF/qvTKRkY5nqAIEM/E4b6IEbAq710E9dqLZtYwwiZ7CShnjGo6Cm2vCkSP8/XiYESaEWyv0O
F7KaE1frUC88dSt8RR1OmeZ91gDBSp7R/PhVh1X4tHqm6gsM6lXJHBxtKN9iS0EdNTZ2gThsWOsQ
/MRkPZZjMV2Zw5K/kPmyP8kYLgz+006WZSIqJyrbRMoT9ITiru8hE13hLMmaLxzHWUqzZWG+nnE3
gLVFIfe9anpYcbDLeVRw7whDA+wC9Pn/FhydqsDiACVaYDriJH8udL96zPeygrQiAWUlHeHLYrfl
gc1bh4ATG0iWm1CeedDLFWBv0+CVLEqKg7W//ZW/w6qoryMjY7rAhJu5dd7uUZwKLWTtVS33Xe82
k4/NGnhYHwMFJ0avnF3znJ1TATfn/i+3fIKqu9o+ypMhRdw7c9Kg50f6Iw9/xs80KOyWBcmMu8/h
ZU6wn1fZimv4siJ+n4gOcW2ReCuLSmtKmjYXk85n8R90VavWsotT8hU19TW1Qvt5/+7wb6SuhRYg
SD7eQbFSa7mLDgbPxZQT/qJ1oJ3yyaZ3oTXXBVql/BQTvUZqqmU6eehVAxXEEuXCyMtpTPAPRFHR
YrcHhxIQVp0zLFAvwULN6jHyuYhefPd5tv/E4QYVeVy7EDwX4reKWnLDOhcfRh/aqnL/Bju1lMao
ndMJCKlYFdc7U0du+dbnWSHl+arqnke+9Dt5t52MvhDiKYZsvgXAoXp8Lw8NuYTImRo2gIz0GJ2K
rAYjJ6YuyuC3O6Y79eNy1bQX3ihA8Q9d535mJe9DQUEvyEOtSyx7URPshqtuvKCdqw3eYO5FV31+
x1UOFq9BK5mtOJtPXIAN8+zY6+5HInVDwJrlb3n4FlbQYS/t0oqRPjVjgeenRVBDNjOXQlI+nLxp
VDCZNVEa4f16JujP71EEOdhKlWIL0XqCQNFDJnNG725IV7UnhHnrTeZqSVly4fN8D/yK8u6sAr5Y
6UNO5zK7yMAFkeGC5EKHbTM7uHYrgPvD4SD3nqj50O7JX7p45uankcp3Icnf59LCOyoAfeuCHEAu
1qngPk6kAOlZvtXICQqor7WcjchOLXslSzV4i410KbP0fd5EHotMEnMFVVPuJtjNLSbxGOOGV/nG
sWWtBNGlzGI3tV1YHw+lUuzjI+ld4++cbBxN2hsXaaFjrqhZnrfiJyNOsgMAsDrGvWAB4wY5EKJt
bg0DP4EhD+83nR1Pk65lK0nXG1bL9iiI4hW+g3nsQrtNY+hWTu+QoGtFXHb8oqq2xjkmTgaTz9x7
+VUeuDcfk4gPQuY2y2sI5WPTSF7iJ5ZSgGuybSiWkBMRndW6iH0Q0doTc/enkbMdqh6IKkbE5qws
mkXrB8BqL9StUQphbT6htvp8ZbweZTKt/B7zbC3oys6SsKqUGBlzBbZ4nNE7u2YIxDhxNCtSkL8H
oFkoOPs/we8qIbqS1tpBQ1rf41xc6QZAGFZDjNpRimhGyNpzcONmOB5C4LfM0GTswshaa+oM/nes
WiJ91/ppNSapJKKk96pFEyOfGHyWlahFd18CLKbv1bEqG+lchqxZW2r3awREafmdUPSxeAPGmJLA
OtZ5gmMK6WXySJl/8ymBx0lsZYwIzJSOhYHEiv2ivXv4Zy7YW7o7l6qGTRebqMiX3lI2XCHhtkDE
nbjpJXNyLwVUindAbmBMoPFBhu87FW08aQDU4+9259dGwaVTwOXgciNFfSWqkBWkVh6dxObzutY6
hv+fk5PcwculqxcjPrxC7De7dmg8Aluro6JXyG2ESSJC3A00IkfTw4Z3pC8nAAn6JrfMbetHe9ty
LrlyiSGxCdwVf46Rz9MBg6CvGUi460e8hhwZvkyqNQTOxvBZyanyBt809xC7vzPv1rydRLPuEmD0
/6qsIS8ijxE0FyR3Tto9/9rT8ntVb8vB+hjQPbrq0YQKTJMBARpGD5udhwQoDdQ9iy3HFQidjJKm
4aSELP1kyGtV5g480T/f+cblwV8lquQ+ApFpDiJKpyKxJgQULTBgi0qNXHiVtG9fLyFatCKDt+Kq
433eSSFN//x09Rv0SyUp5EYqUxxjXE1qBr6BZkevLrq2H2uCyh90Q9CZAk0llSj2/ik1YoO5pz4e
IgzeEulPFSDdMI0HyMMSMb+C6t3/wQFDaGJV/FHyPF6IzsIEokUkBYIENBGKfo/ZeRAizRdCQG0N
dR6mHEhOeiZT8DHH+VWyxweudaluIfl5wwve0NvSPB9Q/v4mVUQ7hKA8qDn4+zCCESrlzO1dDoi6
JJ4ZnQtaf6bLjODbdbumE8faiB8onhh7jFo70nrYxVhBvmNbYWIZrnGR2wDmJ/+L3dw93ZVgf2Xc
25LzPct8w6CrDRcnGzoA+QHLTaZiMcitKjNC0ilQWYuJfXhLDY9KnM7z7GySLZRs5xv/XmuvSUzs
J2Tjx7GTr4M74NyvICZX+y7EH8SUXA1PU+eu3UNBo37U9WGAIHdEOv+oUgagtfIc7TJaaHdVvtSt
MYVgz6gFmXHwClLR4dMhPhdmP0uID+emcNfYDR1iMnkx0VvtTncbB26thNVjmrsjfwSJxFzpOaxi
iUpUv2Ri99czxVvjBCXPpvRi8yY1IE4OmU+9L90wwVpWzZIUrMWf613zqBcljbKIrDXJHBWkIHIH
qWUPG2cuwc97NAs2vEv4JZ9SwOutKeN5W6hHxOGI0c+I3DFpQNTaHxeDQOpbgj0sqktU9c/AQhp4
UHIJzZIfKmbxh/ArSRAcO8i/0LL+99tQ1HhkwMf5i4Skut0JVC7GzVxQCE0F6iDVJEfztkLIUnjm
sFpP/JkIi+2gmRHuMpOe6nfdyCD0nfXRTi9WgJy3iJFowqYUuffr4icvMEZ1Fl2cj9+WhUEBuk9Y
msbDUm3fCIauDi9YGAO9nxZErocEK4nf9W9c9JQkWks8lxSK3IOCac/h92Xu39PIrhyGMK5J7OcF
0zmSgso/mJ7x6woUSYUVsBK6Z/W/IeNYZnkpTChImG++9mrxbbDaY3s4Qjz4reGkYfwOKB8jCqvM
4q8UFAgKEopF5aFohgSS+qwTr4rbowg3pXhVBl9+O0IecV6s7QQWUTJmbYGniy5gokqeDAbT8jG3
RBca3aech0AwmYDBoZxlqU5Bx7ZNK+k4jtUFUWdr0vc9t9y4tqdjjLlAri0IQfZiUt0Lnru4zVj3
0JR888itjxLHR9kmlBWo6+5ZIyMoiHRjKQb2FXcCtaxd7bpUlbtt2TYOeT/kkrytebXbg07vkqZ2
XZVasfUPVKsR4CljOiQFGTHh8hEvtd1JkFC2bR1N73FyerW54lhEb7lPNReJaG6K7KNSS0y2HCji
+0nmVZxEAy/xDOsSv4S32JugJo/GbWYr+SZvrmUvH4m0nM7of8ZuvcBrd/4Q26u3IhpvI/rFRmp+
9YctUVx6Kik5j/wAwN6i46zguhTpU9X8iKE6/KP5AhGgjq6zHleCInm47YvGWIEpHSenDvXMKbnQ
K+YYDJ3RrXEKWowcSO9o7/TrubbxjtD8ilT2EyKzH+RK3h9IUYPpAnw6EZXNyszHHgllCXz1JVWO
RefB5bnsGR5epCsRfEdmwzJV95xT0W0/PS+DhZ5F+yxpcqdZonN+h2OPFyqRJlgtq8R9XF3+Yt6O
bZCKAiFiSy83dpa2fs2/Ud0vfyGNK40ybn8DPiFpwKz4tSmAcNVhlhK8mLAtUHa07uev0s2jo+cS
5jMIZmhbV8/4kLv1KICci5qv69lk24epVaThpoZcaWPQuleFXuMseEFKsGGzf3wKauBDCKSrTkab
eALS3AxERo9OHW/YHRpPgmO+zJJTwQUk1C+S7Ze5qMLi27xVjDoant/PPipmm/ZQevu91kGn16t6
zuUuY9M1F84mV/PPhG3aYFIaAvLwmB/xSD5ZJ+e8lDk08xZrWMxx2VqBpEz2jNukj799fHShHRPN
+n5JnDHQ0Cq/iiBtOTsbmVZ/hJLFxsgYVYAb0ZIG7Rgc/OLAzjrtBqbL8+FKxOYKumuXO2mH4lHI
dxIfzC7jX6vx2RX3H2x5gfm0Bk1VjksxB684mSgjZEPm0ek/NkGjWPbl2FNqjVOwjejYDGoqS0LH
ldfxeLe3MM94fPggdWEwCj5sDJd/rvaPKQjbHdQZiT4n0C7UA4we245e8eK0g/oo8QfzB55Xo7UH
sQAuNK8/vrQaab1vNoTnQnkLxBn3NqHUIhOGVRNvaToPr9GoXyWByxNvLVgPMi2vbq1o3lwn41Zm
oH3g2JPA/3tmJM0ZBjuSDrz9GApJrmPuVZD4/CyWC/cgJ4SewWG+E4NizUt7tYoP1zGsWewlAi+o
Jc0KD9UhR7XH7bilsp9XR6Jxj0hZ3h1Msm3g+fkqEBPJg/joRnRSDEMFdeb5vQ2QeUUvN5Q2a5ks
Ro2iQIPz+z6jRm1nk1DeOi0vSuyGKAPhAc980/5qirL98ZBIH8I1EqaxH9Mcb96vlyMUOjkT3w+p
uAr9E3dOrt/xA4Uq0BZACNnU5tjxEJCTtPeDsiZhjXqYjxXRzx+q3KTpD0bFD1skXIIJ5z54zxY4
B2XkbMj3NoOooYRX5XKPcFTwPTkJd2tJbb5s9YqYSmM2kNzF5oEFxZmta8WeeQw1zKt5GFcIbEsX
eWC2Q1WWOD1qXuZJSqdOmBUJ3MuXuRvKshOEPKhQZn0ZuahxyeAyOinjsS4TAH0Sc5Ln2H0FFK3Q
rXXN/hYx0sipwdIYbq1V+eywXn2aK9keo4pJ/i0+iVdTfA0pyaLFlzzFG430XXnNMceEyuLpZcUy
PZW3PnhwgMwYD4iavjPNgimEvH9t4SCYkGmycUTzoyMJjgK7Ia7eel5v6pvo/WdPzYCgTc+RlVyz
FAgpUPkXIYGj/F3stA5nFoFo9ZBlmp5omOx2hGDWojrO3wr4XY5N+vfPt8UT8SaWwkPQLb0xUfjp
uB4h+lyj7R+r4wDSzsb94ONKvGOQeYeb9a/zXjGBCivDowMQ9tUoDiXi6UBWjkc7F2FN7Fb6fEs8
6JVjcU9ijqus+FjI5iWEYpmZ1QQ5HXuJNHYN2b0azsfSc1M0qgbCKWsiyBcWz/8h3IPcktoJHHz3
M5oC7/oaejEW8jgtn+MT23T20SR7vRTsuEOiRFlSuXZkTlLBoInYeuf0frzWXbW9UBw9JL9qfyQ9
TsNbyymtLtif0sVV25m0ZsQz2Ykxf2i621HxcmKda50mNWXv4kk7M/8XYcB6KJc7OTMVdPvMz99n
jmJmUC1BRZmShmwzZgxNHwyuCHN+8UkJ/70IZRXkIxCYL3hkjDGzPaiQQVfZulLQ1nFq2G+vs1rG
3mkaEmLtlS6N9o1w/b5XSotudpp4ggOO+RgxIlto91VeHLofNsWNM3svpXaKMwI1lV152HAZ2mXo
gjjVAdN86RYlTiVnO4vQiBK6wmTAs6P3IOOtZIRwdKkFQPgEvVhkqNzj7uOxQ84Efwdir+TOMfsp
mFONUjd6lXAOEiuYRzbFgfrbk2z2dPBStMq40Vwe9reL2RCFWI6hkirHDejoSzN6EaQrspWTw5RY
SfsXLO6ez0pbKiR+ujS+PIIOfybt83AnS4X81QQLXSaUmTBwxkQvP70iSsg5xCqHUAQEANNuKP0E
q4pQ4NHPg6eSX/2IKhXc1I67i/D/k9pzqE4e2UBxTtPFpeVmEEm88A7/P4Ci+EW3Le2Nwi4kPat8
uD9xHq+FJI4FO8eVehdq5G6pZ+S3owk15oEL9XbxBX7TUE+xS2dNG5HOKMAWbYVxh/w3AHfip3yj
UpHgmymV0JvIAO5oHeexoUf+hVpTPHp2Eu6NQj1+SzchSIYDqSDySIhr7dMJpWVMhxX1InfecnNS
gVDxcs2lrE6lXb0q8gTmywAcPXmXXC2JL/cMW0YvEi09erjLtkzyp/2lq5sk6bRldD/htXRusuEh
8HDcfvom5ZSIfiVt0xiIes5hdz9mn9yciuXyZGEffe79MC5UUcI4WRSHyHs7hPl5S0vBfu8DL8VU
pHGj6abphkf21cqwArvmmPAse5EAfDcCFyue+KTm6lGci0Jw/XW/AyUFibuHQaN0tbYH1UNm+4q3
+v5S2s/6qPgkerlaY74RMbcNJaGX7RlJlzhO9hA28owptJKefcv+QlPyj4nPR9PHbdIVu4ufcp2i
Cs3ICv/Cd4QT0eNzNAcEfDTjeC9GnEyJxQSgtzjdGrW7DsY5gjLN1vnv2fpYzxMYP9jmIpqR/bxQ
GM0ygnqDSe8nBbPpvH++1aW2qvf2gAzAVAOkFSj0R08b9V2PYjr21QRr7jb+rXvOC9QI5o7NNpXs
aRNB+7UaGGqQG24S79v5VJ4PAcBiQFJGsX50FyW+GG1gWdEXynwf9JV6VkSUHB4MAcfIZ/ROsokM
nGnRlD8CJNB97kRQHnUQESoj6zaw+FDOaIgLmwD5ZfuVL8XWlC342S24G/E07IO0//jt+KYsaOhL
a9o/g1FTFVT2v+Nb9jnoYlN7t5Nzr9qWxR3vQqtPP0er3tsKjz4E1SPADT+FlVHipUPWbP+rl5J5
CR/DaumzVz/5pBvuZvZ6e3kEHkFVzLyNmpq4L6ilP9Eboj44kwVPS1MQvHjZexzZRk0gC20ZYGIZ
4zbzlBiqkSYEztA6QCbXVMvYBVqgunU+mYFU/zIGsne0Nbi9IaiLf07Ktvv/9845sDAangQqq4Ck
OB1FHIsOSv5sYng/ex7ujvKTGEPOtekDukSnbmQfIx6jxttQDCTKrm+ERwtBtP5ZDaWyurpxVqNj
q4UFceHLb4FMURZ5lmcE3Y8xm1oknbbQPEedi90WKVFFaN8G4zM3X2+kdP1iNBK/7EV2Rv7kL/p4
WlvngBxYXg0ZfxDa8ggeidm6+aYuAVDNhPQHg5iy6Crhcz9l8Q9FS96M7xAVRNsMhqe3uaeI3snr
97ILGoUlZ+MJDguZ/2xxioR4aDgnqrXJEW2JVC2rC3MBXVFhAwqn0LxF2xGEXJOAeUaWeVOBVZBz
kh5poBRuIM7nOuL5KAP2sR8cmRXpW7FIM9VfmzaJk5guJu/s8w0Ex+8/jKhkrLt4CV26tcqOXud5
zskeLp3xGjGWqFdJXoNBdSrU/Ng9fVBTOK+Tf6ejSknKh53Em+vrrBcxZ2JEMZPnHeypbG/Rlr3t
mBBgJbIbPG6sgp6SvdBrvFNy4VmwuTJXWXWaKCW/WDzRM/HHCwdDZ4gKHR37FEHTW6ArEgP7/mhL
/JRmWBQDlA5XOtzPGhrGf4QLqzgO3rCkDcDKVoKYPp8NaQq625pdWvlLxpjCsoTp422YOP6dszms
m2carK8Tz1D7mtuZaWmbR1DxWwt8ihGXi8eY9ZwY/Q/+nZf+xcY4agf9EBpREWkiq0iMAmpT3nJo
nWKR3XXOmtUOnxI8C1cyB3iIJMWMY5DNJO2yhDO5pKWPVRr5++2Z27eOETBsmQwgGGsgndDmEsVB
YbecGO60M5pJ0Uwg0HTBdKLCqmZ8RTTTwW4O4PTdfmrsycIb2WmiW5Z9DdoYTKTPMuAwplIkOlLP
unQ3aG0gOdsIx5fn0cGbH3v8/BJ6ylOZU00fqWsvBpf/MDTmUPQvmGIV1clsJX+5XDQzeUTffgXy
wbCDilE4cUE1nQlr8vuIhL9KI6O5CWMgqat93EPsLcK+y6oD0MBCcWkchrXXc800Y+YZKAZ+RfgL
AgBrm8GvRIQCokF9ZIvDSnFZ7NRuM7f038mR/cStkLYE+GPNaVcrHkIyniECvA9+LrP9+VIK9lV8
mWqzao55RaTqkMZrCOk6vKH9k5pwDmdYDOdHV8TDARLH42/lxO0S1lP0p1HJncxfgux/qrmQ3Whf
6VzVfj/nwPgQVBbn0rwGLFcfoyPoqN2wYEg52OKbF3sYwFOX3smwP8WqBSDMuXgZpya4EoCxNrru
/7hHP4+EqCgKTJra33ZirfbmG7DSziAdV1MOAbOaPU+eiiXIotq+BKav9xCWjuoUXrNLlXy6yq1d
O//5odoL8xDMPUZDkEZ/L/tAz8kQv8JJ/0l4RYNdBhXOWzgCC3i//+VV/aRC2StWgjgvIOqVzfZS
qrI+hUP6HxEQi+CTgdNCizXub7tPl+66yQUVqs0uBvmi3W/HCl5+u/s/9H16hYAxj0wI6pRvkt8X
3+NDecb8KuIFreTtuihS+14akXxT529apBsn6u/ZPqK7xyrJVeSdZj0TCYIX01bBor36DcQvg588
vfVkuSMY/XY7Lb95kpouyY4SeuJiQWF+aHs7SUiVDAuhI503cPeREloecNYVo1zWW3v0tEmHVOix
jd2pAcZYSJVlxy4ArD5Jwl7oGhepmngZ2IaRFO3Qkzcd7qcqrHkie6nPVLTu+xG8QJv56/l4gE9s
i3LW26Z6zVX/QL2BuaWkd+tfLw2+o3wUzw2zvl2oXP39I+kXVJyNyStzh+AA7aB691d8MDki2Jxp
AQNvyKh6Q+11P4H9M18JT/DlEl55QfzAMmnZ48Fjjd9APDWzBMjLAYfoN1IJxnc52hwaWs8ITlZa
Y3Xf281E+vV+6HmS2A2RAQ8LtpEHktSC3da0wfWI5exl4bahh5BAla9iVTClAZnJXWMDyXgABUMm
KJ8dRMGcwi+2OlbSwYOv26rqY7RD2I82nFJzfgNzvqo+2CE+PErNA4bOyRBVcbRQx7+ed4jLWx1t
CGHX7whxo7bNmeO9Kfj88n/tJ3gQTFnnFvMo7+ZDrDqX1/oIw7OtSe5nV9TzbGQXxHFiA8rMSaSW
t3klMo2ai90IYsR7JWVBNUiZOxYgTidbbWtTn86Jp4+e2KnJVqyvRdvUMIxUvB20X1L6zVx98zBe
ybFaBW4VE7W3HnUBp8ibpoHuMi+Z54S3nr7PtKR2tLv7ECwPFYGvTvsHX4AzeC31r7j1gqaztfEa
7nyQoAzjHRmKsdzNb83jyvWS7PkWluYeAkLyZJUpKqzwQIEto7/VQ/WJiOlh1jrSa9laRnrV2Ctz
DUEn1RBJ5FWwoh4iZ8eJxPtZf0dKox4dALPo3braUooy3oVL3C7Ao1WRnR1QWvjd2TPgqbAvivmz
vu648osRNafCb77yu4Bjd8K9Drj1gaJzHS85U+4cNSSXgEj/xXfcO5OAAuWxoB1peiKzPaVJ5MPd
D/2TK0FSLNGXheEFUWJlMqfdUj1cn+EkSQZ+4NCd/nZzwP2Chtp+0CnY7G3nID8r7IA3LQBwNi5z
og0B77YXz31pPxoILud6hv4ffz8dahU7HqotJhtZu1XyV4evxLSTdaXfoN30oPO7MrQgyRcSLZ6k
8PbPzjFxn+f8HgZaQyLriPLw4efbJXKG/JvRNlq6YPaTM3jkyPsGcTstK1c9k9LxPk0RyjVczKQw
OXzJyAH9U25SW+TRjqxIQHca5ZuJtN6E3l7rtGrQVqF5ZJ+NIEu8J6yaBmu7eh1I5arH87+L6Ngp
UKg4h7OVZDdDYC5Gu6YOM1j8X6EZ6HcdTFReMlCSouDV29f2/OcwwJS6kjovlVKBe924hgxX8awY
7q2cXNQjQQMPvvVD1mVDe85gqnxbne3a/K5mgp5sYW0Ap7bFiJ/58QdDGq9tAv4jcy5Lokygb6Vs
SNlsrcaNzkee2CSL1g5cuHp280kpIqwG+VGaS39RZKzGOB09+dK4UZ1SWY5z1nzjck2tV6i/2nyH
FpzmS0bw47Op1E1thTmxwa+2G9PPfnzGRU/LzPXuTQpy2ytUom1pkoA8sgE65NvdLrUmf9n3OBVC
KcapXBemNhqmjPtuxDLOGb0pTjIK77HWAdUltEE7Rl+jcraQ8/a61j5xv0gEkh9AplZ7+l1iiHKG
NruufGOoZJRjh5YcWGENhujYZEXqZ7++th9p8iAgHCWRHY9LkzcbhCi3vqa2v66Lf/b+0kiwksKF
844q9K1ClXJWmCyaHbkbOY0hFvgPIWVKKwAp5yRk5dsGKsl/OE3rge64k5wYtQhlnWoUW3i8TZq0
fWPmCEsiB0gO0B3MW8g90o68EZXt8qFyAcjTQN7Kd5kbOD1y9o2P9iwdLkesSqEZYozNgkj3ePqi
7L++N5knAbDKPdEoz6CDcDq0oVwWIoUdPCL/D378Qcgk2YFE+C7RXpEJ9sjDT+kot+NEdg11PL7l
/Xt25sHFsXOKSWSKcK1VikVLOqsZbJs5i8WCVZ0mJJ9oAQYIyJNVkKDD7tYzmfdDFEoqnXIXrV81
Xkr8HEIc2o8g+3+Uf5ubody/lZl6T1g6EqGA8GxQwy+OH/H/hvXxZdZ/9Ba8WiK8D+YH76mKGW9d
I2P7fg0Z5mCEHGdHDM3HpolLjuph2H5GfLyQQ6Ezk0sosj0cTwzHCJCUtuOvlU/OfdOMO3EW2iWm
X8eksHfS96uGbuxtJz/ZM4pqbSpxTRTgkFiDh+pEWNl97eyIF08vArEU3QVjLBeTOGvKon4ZIpgu
Ktxc1kRMOW3+/UkWww7xbAWZTqG3Pgxw9X8W8Mr0Db7uEbx8lC8/alOaczp1x7+f/QSYOk6H2Upi
leagZ3/9kk/JLKSQ+Xu3OBA3+M1N3e8uV0BXfaevSMIMGXft2brroqanAxT0RPxTGexULeYNohzJ
LYGs5Fi/EIpqUwRv7YeWdTks+CMtf/a8uIyrNYvW03n+j6wDboPsXMc+oeqgvfqomGuffRb3PA56
e+zuwu8pf+7zTTg+FRX3kQM7prqtOezMCfrxBlvcCDtQ7Rgv6bn2zyj2LgwebXOlkaajC5/JIul0
e4efjyF8vmXd1JPeAhpj3vl0qaSFxvoTSEsXQuZb9dcIhXRPgwEC8Ei0YE46/ezqAn/p06Vp0tFb
nPu9IyxgN9aAVWRRrrpeOHsMaiK8+cunR1lDHTs8+ghvv7oczcgr/lUWE+oF2xtz+MFK8GJsXj15
2cQpxvqaqvkxYuEgDLPU2NOvY2JMkrz/6a3gSVXLd8rLxkyend3hCZv4XkGOebEo0mF4sbggbsRo
0J1kTmn3wgKOhs6UQS3MN9V4Hn+3Bq2Ney5fBtcodRwpGoQAF1eWdX0ZLWXvFpce82Gd1ECTQkQa
7paVrri6UdCVHl+4cf7bhXzhw+IvGeyn3jKM7Rlnt53giLcb/RWkHy3slIQ0QwQxJLaA4kyVq113
rmtYmNwlSJUKf6niGhSxkwe1bj4V1j6VX6DJ/9b5NqFiVJ7yjp5n9KuDDQcX7WSS7lzN0g3qUJ/y
p27Z1n87UVvUTe/jVBlM8E9YsC0KhGmIRXkPnD8ZfOd3RDaNEQpYKijixTMR62KNgC5lgZFp3UP1
SAQ3zYVvMskUe8Ez8/z7S+P7V4nR6203xZuLPC28N0gYmbsPUEIRsdKFO2gBuw/MVl8g1jHFpVG0
vCCbF7H+jOfppHUZITXaJ5rmuF2EbOHU40Oy+te1FBHW5VCIY48YRjpuq8ZXBZAwXqCXw154MRn0
h+4d8lAYc59OMEK4HC5H2m7jLy3OfdqAtmgO9kLhd1/oxIABaRGqVnWBIEJ5vBoCNu8kJl6onFLe
r07+Ru/tz8XRMZu7kSF+e+OJhPalDHqNMggxFHon2X7XpgD4ec203+Eca39UG1FS15dmytwO6KhT
VGrsoOG4m8CqcQbmbwADSLtfGktd5r0pP2UyH+2PB/myfWhQ+fY/+2niKJkClfqcWDfORTer2oM6
e6II7ozQS318HJ4N7MjNFHQMJXmw6ztdtDWMeDZuZetkPuy28jnnEuJnPICeHiwSQF93sg0+N8UE
vaMCQDpBF3UP1jWnQAaWQEDNZJVVFof7f5N78Ysxyym7VLmnMGQCBN8mgaYQSO9kmBHsfJi/TB9b
egHAZPSKWO0uFEwtJojMdDIPMnMLOJU4Qlvtl+emeHFMp6VJyw6b7/Z13GzVPyvhDtMF6E5OlyO2
d8rdJ5RJLN7AHjuA0UB8/AKV1JBQllRmPeJL0DGg6/UBPq0hA78TwdFrUNNufve9mcYCfQFPLSns
G0u4YqhuJmMsN5/1ZRJNXdlkFOh+xV+RT7Zl4iqg2FFblCTEcL6fvfg7rTkZfWKb32pAfPFqsbU4
kIA0/LsNPgM7Vd0BOmjNGVpXe1u6tRXcsR/UzCKFTMTt356Cq2JMKbJtUrrGnCNNFjs1thRbtMcs
vdH6j7ts4zpboEQKE8Ci9G2SYTm4zzRwbEz6IOWQZ7XyGL/vldzoKyxu9Jkn+cg5x11H8ekqFXJu
CStaXN+oMfk6zsyOgNlm4V+ZysYljrmEyJzglpXrm0H1RXytDbLEmVIZ+zcX5yb8Qb/r2Zx/qyBi
aK9X4ea/hWEelmZoy1nviRxPdU9kwUZfjlbemwZnqixX+kVE/P+W1oR7noB7u7ARE12BSCh9SJRB
snkaz8Z/dbZjvLDEIgjb62dvn/Sj5RK4A3G3NDNQK7/o6REwChAnJziHKvc/bcyqLO50rNqcDrwz
5k0/dF+R2fM6j/2EPYCKWzS3eCr21C0dICpua+FhCIi5Lfz+FPi6dhgeXLc74Bqe6yDqaCUkbRZB
q+jIAYEfza424HxbkLxPiET8iTaXTEibit30apPDKIJ3xzYPUlvBv/O3ow03+hr858qsd/ZB8OHO
pIXI6CWBMwaijnYoPsz5yezHmp28GPj51Zx6xE+ZDEJVhu4OF4yuWwaF0uh9gGOFEIpy4bwBLnPr
Ungo8lcEGsDx3VHkGrQ3ZgP7LLcToqUTBfiwQxOyGB+rYHL71I7NlYdwrptLPbb3Gh6TaaBk2pbY
7LMIsUJeqjgevLoVBn+a9dX8AD0cCEBgkvNCJ/6vR+BTM3PMPdOw9GUAvLUtjol2ptXq3ECGH5Lc
bBY0gjU87CSDmUV6wjlkibY+ZRzsapUdKouHux0UHkVXnviP4WnYlH3h/VdTJf/ah5HClc+MHeDP
R42/qtbZ2dCNKiRWdRqnZyMc64/XIyXCziu9G7eocJlGgbYQS2eiyvY/UQcGnCU7hw1+Ra1BIrdo
RHsKTClG0fSf5bQ+byFMRIijAqE6UCaji+ILexOcccpuErI8FKp3lay+GbE/TYPUqPm9UCK/gG3K
udkt8WhVX22J4S0Y6pQ0py1yg8w2PIlYyw9nou0UuOZ/U+vEhYIZ8KOmr6Cv6Lbe0IjWhzjKvCsF
I685LbE87+Ys50mHfGnKBQUUmQYqxHWSeEx4wjJg9KWtoROOsOp2/A8oNvYSOo73IDBF17Rhyhjz
BFA/l72a3aSe1AwquX6sN5aUoBYtkQ7rlpc5e8UDfLcuG7wI9NDaPuo4JNv/9AWnTKmdZoHsJrDT
Bd3WmenTwyjNE+g6Yhbi1Q3GY887HyADe+9dhamIPpaCDXiycA5ip0naMcf1BoX2p+JfXqMG8aT+
UIBB6sMmsT7t+wNl2la65MfOUaeH5l2QnKUxbs/zROWvZzKFHrJ74oHQyfpkuvgROI+Ebv0z0liw
6r3MBsiS+i4Apzh6e/Lgjo0GAlpkz8pdlzVL5qrC9sfnigPCYUkpiBlsvERLM5u0JYrBMXjSvaSq
gqXpxGqXBqnQLRM0wJvoS+L9g7i7eZJjpTCPskLh3+K1cnXdPYzulGD2w7TUBYRiZMHiN9LxV7id
1Xy6U8Upl6/P9G1fJr6BfLtRGHzLxAAXHAV+tuq4CxnArXG89T1o3yhXsZ0C7j0y4B01Fuot5I0i
m4iNiiwuB7S38MOPZLaU7YWkMqLrzWX2C1YrCtHpWTEB5PT62+bQpxVRvmTDpjryoRQj8nTOQsS2
AHnTwlranGn4YwSJgy0zPve1VIFpK/qxzQzzNNDQcLn/usNZ+14HdT5+OxPIyA5e3RvaI7exuYsU
5rICYPmol7ofn35V3IuFecYIzbwKJKxMc0W2zNi0AKeDVUxKlXjuw2F/QIZm/nj3Ykow+BI20Hss
JoHU7s5T/o3+TCJmrGnL50RNZ+SyY4ff4tbf1IHXwYPzYOoS+HsqF/Dt9Jg96R4GG7pFfeTGI4mo
zL9IzwbxAEyYMSQi/sI+Jz2AVcdgVru3fgdYZl3H4Ce2Vds+DS9/X9mK5QFjk3pqLV/8XnzxGWCs
t2aRndOKFNZ0pN27QxM2GuSq54ZAMMXe+ccho7RqVDvCYcvBSfFzGBVCY80Y6B+gg05zZfVSx1sB
+xxgP02qEuvp3ip1+dqSwWwmzYplqA5L8tnhB/+K0JKmlsCJK0rE9WsTKP7BPtMrSZR3shiY6wzE
6oVEfYK13gaLy47pSjEd8V73EAIYHrYGU/b48T0cUNxSYC23HAZeNghLlW1LtJvbkyrRsY/jQ2o4
Cu3GhBuhFW27l8fvkD1ciCaUg/As+DK0w6baV7f2bVnOu0IlNTHDgVk7m2J1Bg9AeyiVs2gH8ClM
Gh5DLqwFxzdSW4JLHri8e8cpGGUOR3WBeggzn9uyUqexiwxAkeqeH2OTiFbCfVs8fzwLrmVP6u1c
paEciRC8PAsBP5wgWx2jpP6sb5ZJcsqC+0oIwh1M0bLq8J0csSUwNIKiM20YdhOWpCNnMa8QixPV
wMBXHq0BCH6FbKjoxWXaG22as3gNAIXXdQHs7uulIOHNA61YoubW4YiDFttSuQGZDzDYsHNFYW7d
FChxANm1D70uq4eAGykaAUI06ZZhVp3KSn/Jp1fw7bviS7ppv7zdx3uEqYc1dgQ6jIFOU1AXHwH4
odHqjGGZPvlinWxlNHwzDkl8BDfn2Z3TKq3iUzrJ2VV67VtXzdBjDfQVEd4GhSMISfTzRcHnDqAN
MbvAzeCBHo5oxqJR8UoLNLAFGovY2w2x68aiffTcdoqVAQKMg+ikJNoKPhX0tdJS4YtmgwGTEeOo
xNM2ZTAKM3Jx3w14BKRBwjJ9vk+28myNcUONCWE9Krt+LN1s/yhX3XVBK5zK6g+rZJK+x5PIwNEn
vtQk/Ptrgs+AQnwo126WTvhW8LLUZfORlUUattD0EMjQyDXhJgoAAIhSMzrzEZ+UCbxWy69FYNgB
R/Q/m9EOrig+hDmaGZblHhOMWKcmyttstXx0PPP3JIyADlraFulY2+Ca3Cz0QIGod5XWueJc4mJ0
GKbD/0S0nqS51DScMcP94gsh7Ba+UgjN/o4JV7zJ+V7ChLFzc8Elihx0Ffoh30PWkSo4tthm5x+F
/VlawqgnUpaPTQqjyJ2PrPDKCJcAhf9PHjeeTPpTc1b52bK3GFLZG0HDTkTAh7kqzYnWjeGlYWns
vNV/sfC1TWGeNSxHTo2DfPHd5Zxq8J8m7jVTinf2k6bOP8/oOkZDsekp3uPGYAMgbLBHONoReW7M
VbvZ6zOQLMn2KMgThIgLppEBoJVDXjqSw21/UThhZZfeBnz+bTloYi9CzZSqK/g+fCpSHvKnLcSm
otdhRGDVNVtXpHgPQEh19jNrWEeEQArTnNIcto088lic4cAuCTMf+nM3mE2M7Dao2NtWGfudBuX4
hZfhBOMARvF6/UgJsGrSYQlOjeq3rNps4rF0RHgT8yPgAjBCZLB0pTaZh1+naHFRIQjlYROa8Ach
YjuBzTz4MWVbdldsxEKcqrG1Vv3YidEtpAzOi6nuD0sIa64rzArA7HgSP3L5HLeLmkp52QcVWzPk
K0OOrKAxZ/JltR9WIFB11n2C+mKI1uQjzwAcdJenATg4S64Ee46vvAwHnhgeUXfcsg9iW9VCH2et
KIDY8At6BVEnwrlYEqJdJ1PJiTzxkTQardDHsKVq+auIdUYLw+relp4iXGHc1CihEEjW0AuL1G+5
vlDKv1KcPLDuhiTkJCRpBxRVhYVyjidDkadmj/vTIYDBLKiOsYcVof9QqabrhIPpLBitE5KN2SzW
zBwsnfiN1yqP3imu36u/J6/Rn1+PsQFnZJ+2839RzHogpJaF4/3LiN7lZDt+nwJmZ4Oa8jzu0hS7
lK1pWUEcDMGqpExyqyIFoyYDZ6vyJho2jWII5ce4KjNc/6qVLKlHxNJF6A200y8tkvDWR8ODYpsG
qZu8ViqchBrMjtze5U3BZvMmeMbGOqrxCtkP5rw/4TqrF07h1kHm3EnzNxYXUaf2qWwAmKNo4o21
MxApHqLlz2kiQY0lmTVfNoget1yflIBQG5hh8OxcNwrLXDbF27kJOA+nEt8AoUOfS4y85qD20P8+
GGlLRk0Ll2QnBBxe7YGnhBrib2gjc94OgSfsh9ju55303ZmysE2OEZaDBW4N+5RBseROSWXTJTth
cZa2dr2JF08Coi3A3tk9jxHJ9b5nOGaX30/bKoEf4VsvbRGQPjDczdm5DyyqCyJAUtbKmemcerJK
yEr/iftR/+IL/rvjyQCg8fkWpQbtqJOpXcfyOTeDxjsKows7qBqq6QIjqnLWbzC5rb8iqt602lZC
PmYsK68ynRWqmL44eOFBSJlU7FmP2MwsBXbJBg1M4BuafbYF6CkGKfjcQ7MFFeQajDSwyQvHt4bE
3R9nzHbj+0zX+iy2PNZJIqRTSkGjEWwUnBGqqjbuJHO3wSabxxtu4BlfMVnlWfWZy0wnC0IfXUJN
wU+z867mOGZ4VZJrYMl5pef+v32fpqhhy4mH+HcV+L+IeIoCaxSrVMUQkDAZlYCJnY9/w6rC0nRO
mSi3jYDntEr/PIupLkQ6l7EVDkQismMUY4jl41r639v4PPk/lMFQDh8jzwwi1BFd2nDGG613j3/T
JbOMjeickiKfywXf6OENzB1CvexpdpKBdnNaUf3RctrCoR8sKRT8MRYKpJuxKO+7cZHeRtzTxF3U
1LvbTmtXed4TalsSXrFaElEbdqX0jApgMXN0oHY+S5cHgC0pe44RLLnNQnTN+ZUG94ZEd44VfqeZ
TY6KvIFHfY6dPdQvqUM7psGMXAWKK7ErAiq216Ky/sHH86UvwuM4QaWq5WPOCb7agWw2Lt0LmKJ7
kRRRNn/GPgl5YmU2N+p2129OJGWY1+TXVpZrNSzvbFZBgpJQMg43qmO6ePvfVJN7jMS8qEI0Xn8o
60kC7IVFJ6L4B60XNenPbVRkhux07f9GgEkfp35IGfh6CYvohm54r74AxfV5egWyP3ioKTI5M3TR
9pdx8ja7ywSpiZ9EiW5RxmNRXY+9BwCd829uskPTrLE8167AI8MJvphdx+3Z+gC4B4Cy+hk/mjhx
q88D779GooJPzcid2UQnQswVLzBWGAuxQsQncKOKYhmu56JsUNq/ROqAOShWYYxkcUer+dpy+9p0
7A7sirJ0WUTSvpRfYG1MV88NDLOsRFrZEQKv+rmPZnWrfelIf0LHZEgDPC9n9in6iIdeNWs49p4d
IaHVF6Ci74C5dfjZX+0qXrmmmcW50CEhwh26yuUw0aGCWOTQIIoIGQ4lHhupMB73mjB41diE1YyG
mikStmXrJi2KtJAN1lwlno14NfRQ40PFHHW7KvOC8j2bcQgQejLRh3hHajO1IeE7rNTAyUxOdQLh
rDj8LBTVdFzsbmtsUznbEjriQPG1cH22IhEi2cBJEe8CSq3XFTOwDXG3P4nU7Bx8biKRexJWU0c/
E5CRBq3a5CHOJo+11mJ01mSiYWW2DTJqrnpBaUDu6wIyBMD5aYs9yGRuPc+ECI6s1Nu6TlX5/Dci
ab/grw9rpEGtMUXtMlTnMhCxyQTQyxP8P3ZwXBdIf+RbcVR4Pl08bwSz2+tHHklcSosZ1aLiP+2Q
U/74YQ2Yjai/uJXp0aZd0BLT2VVdVt9bAHe+Ff+Fd8cIPjKZ5h9e9Xii/F3oD8SF5UIvPKhQcXHH
WY2mx/L4NA3oBPEoYehtJoBtxLpATa42+GUFa1iSpKHi7xnMW+q5kbu7QFu3VcNxyAH8pww4WY1N
M166r9m1Ve/shuNGFiEoOtijss5OpGYVVJlrrnAPirXRz5qeJIlg780BCDTqWrztZWt0cQ5+ycYe
dIlYM0S1PC4gJCnwUkvoH88bNoAV6f2LLIXcAXExgUn+Z8febXf3NBm05eo3/1Q+trWz8NokEwbx
Gm6uWE/rP+pFJwbuRchVHQwt1VHVBnlCAajrwbPIvXkExlq0yM0dfT3g2QpUVgp/KUgEeEnqqQ4s
+hZazNNFFh4PYElmydqsF8639eCHyoyJmth7XMWiLI4yrPy8hpTTqw65HX4W0fQrQp9S4VE/jrnR
/dBcM8cGIMMvdtLpRa5oxqcvXEcfNwlNrPw0Sm2jfGGQmphpn/gUFgTHDfvIHLpEvVNXBErKhSAX
egflohCgmo6DT7JaDhkSo/MnypEUIqGVNLHSVugHACUA428ezIFjaxJzzOuJqNwWifNbA1UTisxj
LjlfC9E+4MU1nFuHXiTWYSM8TSexNUjn405u2jNNljD1d+Y1RRfW+jv6lvAf0DJaPaRkXPnZaI+u
RwntxS9CjeJBesJC+IBtvsuNtlUkXSeRIV1ft82/2rr8hNAX8HdlOw8wOHj/tdXZjOkmeKr7gu40
hojPmGKtND1W5gks2VtuFQ700M9N2ZrgsNMRrdVf8rtvS15fUqtzmYOabzcIu/llMumYTLAjDhYM
b/HCn3mKpWBv/CHmY6Ch1D5fDcUx1No2OUijBU415ZZsp/895no68GTjcMhD+SRoMQ6t/jeApWId
awf0CJtiB0HjOfkv38JN3XaiEWqXmkzLC1Y9OKPlIOGVMe5wgTZT3KmAcbkAcTWMtXBtGW1aPivD
RinlVvmqqa7PFzUbDgOwknA8FfHA0n8uotCXyHKTpPtRFmYHWNT74qWAQTfV6xKagNl0+RrWDpr9
TkiS5YH0iie2keBv809QnFTRLc1ZapZLGE9H4HCUk/mnuiyY8xo7u9VH1rhzqte0DQT5z4wLfbeY
xfaVGct44+TWJ65s03kP6NIrLLBz2yNHWoisbL29PnxBSBbjxcPlpUW3yboE3LDlcMJK99U6f5Ou
I3QvtzdYKxHpShKF4SJE8y0TJKZX/wTYJgxl5IbAN6IsiwQp45BEwPE3OgTHO6KbMbfOokb6ngSb
xp154PGIEZkXSGE6QId3cCxkD2bIeTrz02a2eaDkK1Dbmc5AMVDr6/KIB/jd9KkM2Pd5tuQHM6bX
ilhrqUm2bGCO2KH6CvNiPAI1LnFKCfOJvKD8ZiUjQUsVoRcIA/kjaFRg1+Yv18EjKOufZX70FBfZ
NmGui/7PUYcIPIv3A96BAt5sJR1gzRbw8i+xJGh7kdvbPB4KY/JNgW9AKPwfpkJetQTPkShfv27V
Hn7Cy6i3JjXDdhGJkTI6JcIKjbt9nMDUe3Qb1trdp6ezlsXIKDMCIHHZQW01IpEWzwYQMsezOWv2
t5Sfh0qj2wGMOPYMmCSAFPrjvDqns4e01XCTz3p78NJahrusl5JVsiUqlgSsVQpbHoPPWdTZEsPm
thbgTW7390mnTv9PcpU7Z014khvMKrHc4YY+HR0LY4lbE559QNXGYgXxSVOOVX7WfXHcnxr5Xplk
hCGoyUcy2ZsaWM/MT72dLmor64LoTiDFJBPyBQbZG26wLMATmSGAaDd6UPkgWEErtxcAbBoFCnmI
nuJo7YGuyRL2BLnWDN6tHEeTzouMWUwo7HuBiD/r0x0BgQ+lcH5nWspbbXrJzDcy3KKuwaw9Ctbx
4HVAbZMppbewahor7UnEaoMIcr2LktNYuHS3GdWOIG7oRKS9Xj3q37bCUpNiBHD2n2vtxO+DPJV3
o0e/mfMXr16afdM3OdzXrlrazjqouWowKLaC8YxwaA7/o4/3nVuPSQL7e3fF3dcggJ0iJT30XZSc
rvT7dd/86kMFHfGoTLcwUNy6672M+AQTXKuhdLqtqbTC9hricqpZsuJBkYK9vNMCCpctaB3szTBA
m62BiDDzkR2JQxrKUcY8klS35Eq6Rw0Orv0/GTEAB5iTZ97jaFgREe94mbXcvgLILE01xYpb4r6h
GOWwEf4AzxjSn7HPgYUm36lsDj5JCeBI4kBBUvjX8P1ArNa+R2rHZn7VtH00dYwnPCUXOiHSoRM4
LtHJIpdZ0MV1tnWRy+UdN5N8OISgB5FKnLzFkoJ8c3iSUYTLS+L/ECey5wniQzK9aSJAGMZPB1AY
a3evwtSHPS2KvWgHjLNarZ2/lTerWtUax3r8s0jDIP0DEmZfGupOp8FQEZaON4W4H42BrwM1jErJ
UZAGH8fs3da7eBr7PxpaMMixEnfbhwQHf8QefXj/F1XO9CqlJvCNzM1Ck4Sba5rufahzm0jNvyq4
lg8clm2Ax5WlU+XtlHQDVBe4hBFl3H0XpVZL1dBj1cEB82RWIAZhl/BiCTvzKR8FeM6brh2vd3fQ
5F1ULyUDQe03GAIlg28l7GwZgET8bM18g9oM4pyNIhAA7AryfZaqxKCLKVITKCXTD9WVWX2cufCu
RrQJBLIwvZy+jo4zB9jtenmtK6ZDow/y/PEgnkkrVevPJpivt+XJ421iznjyeSjFCtT2Bs17vBNW
i0M4Bi29sxrhFbHTkR7juxF+FIyDgHRQb3GR0NcrqdhSC/rROmCVQaJUaW0GP2FrG8H6gCRQoC3b
jgI869vV52HGZBSWKY+o4oxl8wJDLTgjFJMT6XNUsu3gAuFACko+mA1cUXLaDkDYNCKo9cfOmoWL
n24swmcGkMo+yuGqv33lOXmlHlRvxy7RJt1P5ut52dn65AT1XCIBU/YDAH9pRexluXF0CHzKYgkM
SxXKvlL1okztd/PH3yaHKeuASu9oXvxORehFszJH0JEYhHIA15pOMT9qgLnRFfd4T0n0ZVT3Frtv
6J5HvrAu5Ly6iE6tmPGsl2VjlKMZYJh2fbAbfTPux7Cn1yMtjGXq6zvwsEkfI2TfKqa9HlqQ+Iik
4rQYiCO7dRBLS+a3j2DhvSc92gFBTAxvdDtEjPiQKN2LreGaWja4KznFB9FfvtinEgcGJn/Mk0D5
VivgCDG2BzoDTghapDmFQKThCnY5lmyDPdQ2bcBeqPOMfITC4NNqI9qt8nHkSvuluzmrIkiXvkv8
1vgIKc1AMXMy+QvqA7vlO8kuchFadFbs43Tauk50aXF2Yh6TyCYKqD0HrkmH1u1CMD2Txw1yj3g5
mwGQhYcWZ8r4htH2qhgJ9HmLmz0Lm+gVtaKy5KjzUQQDhBmO77qbO2n21twr5ixTajzQDbtysAa/
En9aJORZk9Y0opYJxgqQqE4PF1gpcVSAI6WOb+A1e8dA/d1Q1jgBVcILNb5tBOVOFNuhWUr+Z9bR
ye6wXxpQNNvXmcdJxp1aFZzkVjaXLxYM0A/bxg/vfie8bjWZ7k1UFmXFYo4DupuBoaaGC7945PFn
YNe/uNRWc8OBJ8fLkdPPmXSl2T+0/iFdUiOf13dUsZG6ILB3HV9kTqA0OGDKK5XztGS7h425W3iZ
0RLMghhe71Uhv17AP3aWptad/Qawodd1hHooLkcHLAdlEvWW5tOyDBKfXMi4pamlJsoeATtZixFT
TlmQ+XIbBPlgaS5rNx4XKTVd7YyUUrgABo8ZPMMHpyXFGrtYVFPTX+y25jaSyNJEkh067ECzO0TI
dKTUO2Epyal+jNeQyrt+yFHTBtU+pzYfXvfmR47ObwfuRLQ5boh2PGM9PQEkmuoXZNfUqBzpVGXi
6Shx9ss1hdAbhDOzA9JtrRSFY55UNPw5dpnddlwKzN6AKSgocn+GPJui4w6200j0p5iSPapFeRrM
17vETkLofd7DTSFvPooM8jWlqRRbMLSyou0wLYs8yoTLvedxROKgROrYIvTzMTKg0E/A6/HJ08Lf
iyfXSV1LIbyhyyf7LfNeu6lnku9WTBg9G7KbIpts+sKUpF148kL1fHTiopgguVLnuUsRyQtj3zcj
G9YuVGIEZANSicJltA8A+oiNOiVltPKHTC9PRGbLXm+qAHkarX12We7DNrAkkDGbnsVGzixELNh+
W80jkPKTs6xxcsrsHwhGU5VTN0sU9iYsmHt74BCIigwK6CUf93YUAf+oMrACN84iPVJYRNSTZ8Nn
TFCEvTbBdtGTX4I6ebYsL7yM+/g3RDr9/6xh5uAk3gTme4uHJNvElXtX1H8feF7Y5k0TYwc3hDVW
RqbVb/q6EZNhaKLeklS2zAI7xsTkTlU88vlOMjwjQcVg7GUxoKFWFLZWRIBw2GXiQ5lFJotflbMa
lvKosSFlZp3qMqLtAVTJZ+Cb/m94g1XrXvvJRv0Qf0+h1tZNGg861wCVYKB95cJj7cdOaH0xy3Ql
dfDVLrP+Eh0+BhUP0flywiIGNsksOOieNWi6BiU0oKKK6xhuWAiNl5rIyTziWYnJ9f0Y+uCt9tlm
dUJCleL6rkWXbNu+lQstAJtOWxoMZ+kjNjRjNoPkYK9t7T7DVEFDWFi7JasVLNhy2FZZBEMoNc7p
yZIiNs5BxqFeQX36BLRZWV6jd+2n9a+iy9NSV2ifFG7y7BAEqurFSOU1wAw3IFxf2PufpTM+BeAv
7wdw6Go/LIVCTPDviB97MFPiOannxqidWcnGQ6FeZlzYIGCv0hwQQYhxSAKgOP55SCdyplWn9nbl
3HYP5TjYpFd6WF6gaBs1a61m1P4as/MF5XckFbZ0AtlPtES7WEs5kBF0gQtNmB9lRgGlDQIHc4Yy
EzC0ajKAdqnIVbkMDMS0OCX9JR5ciXJ2C+3Mk/Fb06ZK3MyEFR0GckDRUHEzw2b7ao7qaZxNyxHM
bKa2cxdxKX6/A52HEp5bYhcBliVxPgwKOLtAhLr4+4LXuJvGG4nQ4k1iT2iw5FOY0aQa5q8tYl44
sKA841wztz9mt2ayIvlieVHEX6S5XELklVA1LLWNwYdzAPixkaykUO1Q1KWcf+RFG4QM+qM7tF8G
NmyCTu0SqARV9HGCwVB6sHXYjyb41n0AZmnY9verB2L7BdYq1lppGGGh9yE4QIIWMOcgWWHMi7P2
/bAuX0b9AM9joWo7t+3m7vVVFWWdq+YRMgx6vgqenl+gAD44JsKq/vMK12H7s8TqR0l602GNdGFY
VwKVIHRipCBcp0fXIo4y5aozuUZ5sGXwYDDgPbwl5DmxZ6H0VU9Y57rP/npTVBpXou2iwZ1mkFDg
75Y+e1Va/zLeczjRePt8xcb8aRTZyzD0wZUcnuIWumpOH88nV0ojE3bZVC1mJBJ1C3+drRH8dhno
PEWd2Do7FSSu35PMDZkGcnrn7R/BNpXCMwqZyqXeTxiqIsRerqX9Q71/04/dT6PFMIP65HGa75Le
uN+o5juyzsKaIalLdIM4rz30i5m7tiOvVqtgEsVGMw5jwbHrr5a6bhpgs/vlYRX03LoE8RY9CFQP
VYYNnqO2I59oziBSjkRKKBd7x2i785EoyE3TgeDu/tIJIwW7IvzI0T1QLTnj4JYnCSreGExPVxpo
YA4eZFYcfHr6H590D2eqZjNB3CfgzZhLfkgrfr5227b6SYZFRVu9h9CbGkfpQdrn+rbIccy6Nnye
1HQtNsxygqjhumiem59/iRah56gxxxcS1bdCQUt1eI7htbjuEN6dPd1wTGN1pP82Yqfke8oEJzb2
UL+Y3yRXpIwfz6AMKb4KY6EdMUkoYzInkpqR/GLrabIBfFs8prxcp4iLITC//mIMU1aVxtLngw6d
A+mPIQ+KaULbHIad3kdcL+LiqX2vz6PHQOtvvjrtn2012zGVCKvDToWdIx7n105Ap9EQF7ygRCw/
cV23T2Ftwqc7EQ2PeMc6WydX0QVg6CgCecpptrBxFSn3QEd3Dswxz1a3kAdZxDebXS4A65HerkPG
qlXaX0seWH2XdhUr+UfPJah26dL0ZDKCTwmuhje6BCk+shriTmdx+0E2GkgLVLPyGTOaNsi/SOyl
WkI6g80zm8+GtHgCYEGosU5bNlLHJv+tNxw+ukXQl3GggOXqULtvtqH0LBGSxFTrx4ZfEe3HNEJD
K+vNMKdDEGwyWNSseBAvckDcJOvbI3H66SsFXOd+Cp1UkQrt59Kp0oSTHK//knv3tBW+I59UmRQu
GfviGK14P9vPfbiQWKopE4pC5cjAqSvahiqP6UYaD9q0ZTERirDu5AaXfA5tNyt4VsebyL8sZm9E
p5Id9VhNY91Hs75tTdY1rPeqJph/UBgBYfDNWO1m8RZAEaWzqCUJxUm6TagzkGGwmaB1qVV2uaUH
LqBE11vEvB2sjEG1Tx/AXAiDJjM9HPHB0t43pgfHFvOz+qtKXZn/Ve5GxgrBV4yaQN+ulwlGsi5j
6GMKALMYGNC1ArCtqcTidEWPTy7rZ4uFZnDiiPGEw9v+drSyD2SCTSbITpX63rWRJmLhGLBRIEbO
3wVIt1HNGmnNa4rOn52WhM53cWx1s3peA1ACXws2bvcIPSKPfpx/mnrPzvAHF73U84A2f2uOw5Bg
po6BYqTHMyhA9g073coSYvUQw+fYOo2Sf6oHBQELmRVZHKUGJ18W8Ade5w5FK7pVrR0gwWTzVjxV
1TYZ7Ogbkd4nOIT3c2R+fotIhSSm2O4QKEFOGRm32TJBIy6qIbZhNKmIA3O2j1fOziv4F2Aj5tP5
0zsF7YXiCzi8Os+Yiyju9RqaItTKFvJENokG5y8JgBp2qjJTri9lDKuJU97xMUL7TZBRJLQ72kPu
NQTPcHNfZknG+aa8jBbBfB0jNAA5pDIaPUY5FxDCZiE95N3sTR3xD99ycFWM0PPeO+G7zysGmPgT
R6ySBWeHC1bz0nserN54P4CrjJxzHuKuX6Mn35e7Hx3PBT3+++TuWOkbJ3CxXWiJ3pYIL/yQES3N
6vLBajOF56NFtMAwMCXbRvbYjv6hsPNIM/sdYXvgK2PTOjP69LiYT80XWJtfa+G9H5V1zMxrotxu
sptMJQGpd1g+f1zrkEANi7Py3NiTs+o8EcXOwtFxrye276y3El8fOQlXgciYH/aFGl4+rjIuVTpF
+owcbVWg29pySLraHhm40ejw1adBbqxPOb4ZpGIZafkL6eFOcuz48UHlk+gf2j2oCKcDNljRR4td
LBBrVSy1ruD6wpV3F830wVtYHbCvONsHL4XMPPjXaoRWrQRXuG7N8ersL052VSuIa0Pcas3OQjOU
OL85oxFYCld90uViQXNtviQlBaiNnGp0/CAJYmppq8Kfr/RJWpLxDVdV7Cqn6TjOz+cxc4v2snFe
+myJNRieIKdzO1fqxvFQzWLq/XuDmie425HsuH3gSNhktZkqrtFSKCqcycStXiNRDMow3mSQPCLX
DfzLf402KnVWFQmuaKoKpYu3hsbNbZyuO75h/K8IoI9SvAJxM81Fn+1OTXWFm4XyW8LTNhKjo3cG
pK2trRwit8sWvP/qCG0Zk0ETCLe8psv3yCE7f56oSMhXGGgaGZF5iO5TX3h45TVZ83NKzGY6Er+c
l01r7P31t6bGnDekzYtsGpq40vw7j403FAmKfkI+/rz02NXgqD7715qxMYt60UYPpSfCuDBNY3x/
XDw+MwQY3dr62ERsQlIru9c7GxYPUqaeDcnJi+ZbYcgb5zO5mn1HhXbyeuNooZnZq90yt7cfrf5u
FgQW4QkYTuaBzFLEMJUHwQVAW2c47bMwraD7vKiKRMFu1xKyR7XxWwA/z3gH3Tn+ZX0puDNYGxnV
kBr2bygxoZtm4GON0xlVOQLKLBrGtiTOjbsHJZPzS5NRTH5Z6v6z5/C6BlWCncXlm0J5zG7CsQeg
hsXEzvXYp6EdvlTXyUtu/CQn7918Ecm1WTVXi7pfvjjM6OPSjLj3NlJDaVpkYoOM5NsSA1SmiX5z
Kv6QsXnFGEyCBQXbCPBi4iU+2QkjryJNVqA4O+i8SAIegm5q6NaPhR1o5QA1UIS9G4vfPINu4/8R
Areg1gPS5QZZHknerMp52uTjhvCudxnS0XZ9hC7mFIHz1TxBQ6bAE7fnQoWlR0pY/TP0yg95EnwK
ttOt+qknuxeLWJ5phiGmie3mt9H77D9JEA4obDvNgEbx4ceZLWOt5g7jRreDCYKOqNrRvf/3BOak
/GN9q+yttwHd1aS6HlP0hbuGfeyYv2OEYFXTfqZjZzD+mtf9XJOKmv111xAVSucgG1wVHt1EhopJ
lRf5Gqss2Gv3PAekb9t+sY53EBHas7GvjNN7gazsohdnydyfcprKIQA1YJMJtsA7Uhf5jwr/4rW5
k805gZXsUoaN3awSPlCiy59eZl2KmIQiN+fm0GO7n5JGwg1jj085WNoz4qXQUVijM/aAUru8XzRt
VLZY6DjVZE4nO+JI9IxXFFLO9vLjXEy8l0DRXWwOfboZV21Ke9gb62tjIDn9qaspc5nRrEdKCPmF
M3ZEs5D/dqGltyNcLZsXnUeG6wKHvORImT6Mg5izb2crDewlJnQK+3ZrxQuMqP9XnwK/xaMYR2EL
l00b2r3HnUbIMeHB5UzXxhe/mLFcmF0PjXr9V+Ka268aW9DxYNxgdTBeU12yQ7UToHnFVBgzp+01
vXH8mgqkKo4en+u1bleDg7fWkZsj84eJWH/uMzTH26l/lK0ZpZCzHJLteZncluWO1s+rtD7FR7Sv
h+0ont+14RMnBi+0f5eLXUZQub1qCiVLr3HcyIHnJZjs7tl9KEfFMq+ASdyZPbWLfZm4grZQsViL
LXlCj1hd+DL2ai8SrF+IncTvDQXxXNDp5RGv6pgCsaSVKT0Fb6ymDLNk/4D/Nj6FHKjEve2Fp3Fm
uO74IE+eIyLYTQjkDx2Ekx6Lj9G+XtVTVdju6hEFg8h56OBrBoNXXvzJj70RtxzhOVEqrNjNo3sd
ftYGstdXrpG30H83VSLXWaZ5kb6O/yjYarAyKkw3Dg2JWhzRwUsWhDm7uCH+OJLQqtwp0h247281
hW7nEUEohcqCdgSO0aONS7YfTBlRJV0mql+G3eCbVowcShLkGJ2dQxLlYLKrQQl2aefBasUqyIpI
nETq0V6HnfbXviP95ttOyoOdxRRNMzRTS2sSB5ECjHb3UmdtXbU8gu3B7WKKTenoL3JkTBK3f7f1
7qYSJORdKwjki2GZhpx0We099PaX1gV57LISBd7wErHBzb2LN58IYIqVIaPYg2N8vWRWtKVdqwe6
H6LoTbLcLAingI/7ENpDr398hODidc/HfTbMJAiaOn+icgc0qQmO8DRS+umRE6rKux3+Y2pD91Wa
+ap9rTp7lP8EwkDFBJBMpZnXLEb4auHqN7b16nAzJmgbCQtouCBJj/1B3mNTM0G0kneCBtznsiTz
3o6X4momgetwC87UTjhciQ6MD/1TMzXK7PlAb2QeKCl25mWNQwfLuP1v6p4GnBnRZB9xsrz6kfSp
T3cmyRRuZiZ4R0DQ8nW7XoAbvfj1K/Orh/zeEj8N8Z7lnStAkIbekWL/Y7VHIxgEUpwjnlnjnlq/
BjTicsEP/8DfjCdpyQsd/rpk90ahpV53Wza7LLLMhwnxWkAQdrQ2FWYVQyVcRa53kr03t1pxqk7P
D/18AB4RI0x8Y1txDnvetHs8R2CtTVzxTNWpsFIhQkRtdPZztlxZUUGLYSkpX0EamfIpXMltrOJQ
XswsuwR8ytm4TFZHy9IbA58XWmVGtPB98ZLpv51/yRmW5cCk2proAoianilCU3Qt0MA4ueD0Ptbe
Du0xYTcqVjcG7fRgbUTe02pWnh7N5Ktpvhs/O94Dd0DT9N+eqZo0L8VeIWbt2hZWNDwM+17xjdah
8qNVL2H3NWDgQXRY+mGnVyg6Qvp8HhlbxTavUoIOB++VQlbbiXApn47ZzlY6+Kr+kVNgRIW/goWo
tlDLCJVgMVE2y/tB/y4lNREzoP/Es65SULNppFSZEAxL7MzgzUZa3t4Wufpf42SfvWTSYx4zfLT8
7+arGhY66hqdVs1wUDHJ704LEbRJt1s7iui0wSrLB9xJroEtZiDhlLiehZg7P0sZeJNmue8zREBh
NX2AfA7GiC9zeke+oaJsJpffAv5dnHkX3ECMoCoqpVzkmvrNZLBBkVK4EJ/Z4s6XSJ1xabFpJZqa
AQfTYZPuiGed6DDyICnl4+UsM+xXnmgNlGigIgze/QY2iWZKvNlUVNNO8fMZhLovoBCm93bJqQ2N
Bt7qdnrDvSwXBc33BvfYjwpd2nWrQQjL6jcm9ZwHYSqqc5DcsDtoOfah1PAd4RPU0bp9nODs96A2
aVxL8sOVXU3EkpvvOF+t4XUg3xEayoDwpbbGtlFI/wfBryJlQXXXlMfLYdw5eFbbzAOA1IYdXVpE
wB7KCspPsCE0m5AsLqloECePoz7ufgPdF0qcE7h5zOFAw2DV/Ahl1lmMW333Kqh/2Nxx7i1xkwki
4kW05LRiQI5XcR4zVnsvmpLgmfb/ZilYuL2+KnfgAK1u/jPnKRA2sg7vXf+qIIBA73+QDtTAsQkp
YfA4LwCpgfF1NMwW5lGXMGqMPLhTnkb6GBCPeYkPp/CoeAlFt9y/Er74hftE9eFZvRj31/RmE5sS
KqvQkqu7poD925j8mXPy+LFZuoZHnlc4hL5qk0ql72IvCUALs+IONZ+ItJU86VIEgsEiOCFQPkFF
J1shQX1VK2BnIVjfw4m9PrIvU0GF1SHjlvGoU5O8JuQe8c7/qO/LWdFBJ8dc+AWNLNQT7NwrYVTK
wO3Zlej8bKrUur0Bp28iwidYqoq72+9+4fo/o/fiIRw/fqU/VqKIhehwEwB383pF5Vw373woRGph
fnAqvVscnGZVpd7eXzbRUHSmEo73lYDi3hHc5+LBSPnqu79yq/ytEmsSOV5nRRFGWRNvE4aQxVix
pMYXsHH02qdqh3qKdGw0vR+LHCJVst5bl4eTdsn+DVUydziTNoUXNIG28jUTFI2JTBJp2KcjAbqd
zGzJRxgp8hcf7T89kkAZTwmZX1GDEXBbVLtFpgSTxP0T6FUjTs9m1FDfpctFH+ZpU801w++tlw8f
BGr7Fn+hWTFYWuJR3FchRr22AJqZeM04b60uIh5XEK9Qs/PLJj6venbDY6R91IiZlNc3ZtocLi3v
IIDTDfFcWR66JGv44uZoIBi0rywpIQKnAt9GqtoAepFsBsGKl7zGdGx6iuKDLnTh86SP8JUFo/VG
dykOUmxs38K9POMp7uQkzmbXDZrNUCyoUaBSQpj7C0ntWBlCI5yH2DVB9BBIeQiTCvzP68aSUXZ0
dRaFUm63bSHvyf8ngs20j8BULOPC68BO4HuWf+MS1Iu8Z1yFQMXQyhh145ap+6SErcLZzWohMJuk
vp/LoiuoA38kIKtt3E3clijt26an2abDcPfjZquucfIrOyofmo7w/Iu10mGuRzdd9Z3p+IE83AsP
71wv5fQ1HjjozmXYa7Ys2nSqaXfoP5F6IbCag30NZxv8a6Te+bF3l5CG14tFuBYOriFYKOYKWn+h
vselVf/4rYsPZ/3FPkxFRBF3gHpP1Pko9KI3U8u5LM3K9YGOp7jpRswaMTLTx5oj/pEeWYlcw70P
2t5xFDBlVVU0n3pt5r+UUapQor4T1/0k9QmlzayNiJYVvr6JaoWzZ4h1iD5WrH88wsWnJrFswrxX
phIwsEQGHFUYQuDt24YfCpZh/uuCMszx5R+qpMADBYOKSzd2LRxP1FVOBF0ZC0UjzrthXQ9W0+cB
g7xq1XRlW6fda/ilQlWQb9rLLRSAda0a6NQTIhN/wp6wCwoA96vc4XmLwcHjpQX7Cd3hIONWtADi
v5NpoYTJuYRxhCskJ5m5dNiKaCc32E8kNr7op6rSfquypfO0wtmLF6a4fzcUUWJp4gYsqIwlnxX6
kEkvyHdBNAiIKQevmO9R9X7jTmJU7oonhQjQKVQWUnbw/b0mcU/u/8BO5M0RD8rSfk0goztczqjY
uOPpFtULcblaq8/xMkHuXJxTpEUAp7BdoUN+B6VkmKJaZXisixcLZQYAOPZgbZZg02dBK4B7Baws
vhrOiKT3Q30qT1JMSm5/06ZxQXo0Aq02LGWOgfZ+lAhGxjWF/az1LDWTAGHZSWKY21A1gi62Bh9W
XHIFRVy5kXyIozJRbxiU2f36enCSRS8lUeMwvpnSMaOOofbwc0E4cqQuZLVYGjk6xLLmA7XZChnL
3o4Axcz2MDtp3WqkOHGo3sIhcvLltNj5FfIWepVhu7GK87m4G2ox7KHG5bhOTd988JqmJh/nwLMn
dPYZIrEuzr5tuuBzAyhcbzOaTzXYxHdKN2n5z8aDB/0P+XWODuL3BGCbHb94gVkZW8NODW56lLEq
drmsx/QdNSX4RvKVbnQZQLFIiVoii8TqNz//4bvPaa1GRDWi1HADP9T3E3gvXRV6npzNy5dgmV0b
y4ZgUCnVaZIQVLBRXfw8yM5Ole1R1k5+4c7HV/BAOj9fBfxAoxULDalLBjA9AcM2fyLYFpFaJovZ
ONjKE5yPfjhAfX50JsT0POV4laX7WUyrJyaTTziesWW2QQgDe/7Z1g4rExb2TSwYM6ARL/GHPjOv
9q4dwNUo5hU5WgoNYbToK4BucAwqMQw2zPfQhK3zwD1woVdXgsg4KW0/ZWEAAEE12++tsIXcqsCz
E/F/jAOSwdlqfuy4ldPuyESp+9qSqDMT/FfLVLTlgeYWiHQNufXatcZK3Grfj4UNqEGGl5XZvmar
e9blIl/cv0LGw5inQk4QqrqZb4g3c5EeAH6amR74A65m2I4o9NXcjEYw5wfdz5TX182RxlIaVecQ
SrDTFcVzmVCvM1m056bs32QKZF6D38rLNdapulJEPxTo5pI1bBHJspYKMSei5ZGDfAE89gtXZmKv
bp0xh8SpoIUiyE1oSylVD/BppM3woXOm/yLujA09T8OORbcwgCTHuJghVeP+98llPKOSWE5uNqNK
LoucITb2reXsYDKUQkr0iflmxsXPya7Fu57Lg3wR7R6fKl4o4Q6icrZ3jbSgM+xRdBnDc1YjeDml
gBA7mKZwTfrw5Fc2O7lHCFH6yvp8u6csc8hUB1f3NKQOEartKkgjJiCCd59uNiSJJnggvbsoVRY5
zP8K0O8t2+HYtonMR7iLD3qF3gvqdNvRIw+glNyzU061pHK9QLt1xJsYw3VDW3E0IJdM53dNCvTX
+/p5Tfel34UdHmu5zEkr32TO+vDQ7Rug+2Mfz2Mo7UYGRuul5QsIB7AWs8NA2VWAL4XJSi9xzsrZ
KX656ib/47ag89myZyTsXANHHdbEvFsUWkojoXae7GDUAhE9TIVk3iHkveOCBMbHnOzBdfPASxMx
1PKoial9wl5dil0ettWgt5v+g9A8s9M/sfFz8Ru7IQYHs84POJKBKfHlMcmJ/D3+o0Msbbwedlqh
XhqR0TgT5cldy/cvujBOEVmx2Je7fFdfjnZkYGRHnMDcqeZLhIATL4pLqdkMPZMI7hG4QYq8xQfu
dgS1dOF5JE9F43ZHsiWXCj/vXkzhZA+gRb+SYKNEhy3VP8TuetTav9fDzNtb33H0aCRkTsAgnJQx
lcjR4EDSgDEsi0lNW6fz5V/y6J09++C/YBNNskQ2tHwPicd2vghhjLNPAB6+kbP2w+w7+waQqMKg
xRtvSBUESSApBsHkO3TtNwUEPVwsH+wR0eT906DWYL1magGwUq/TZ8kojB8AjuIaFrdsd9g3DExI
rQdzEB5A4vHE7XMlIzQbuzI1b/mTt+EPn4cbpn1PWHRLjbqXvk9BAZArHR5MiITFBp+DqTPsFV9x
efMAZITaUtfQkvhvaw6FuD4p+fDSVNOavwnJF3SEeXseslakLjxZS9jeBvUOYnm+bZl6bp8c6sN/
SlxKuadu9wtJiCkB9/Id0NTelCKgcdLsHjiaiAWBxarNXB1nJaZBkns18Lgc3OEHRUrvrlTHI7H+
0Ddww18uFzoU9r4DS9l3N2c4ue+TjjTBV+fdqII+E59YhXE9A+DJQpTasZ6Q4KT/y7LPzK+B/pmM
wu/T6cCMwdVfyBqc7TBmH09IUgPFjZ/zIARpxrmms80+QJ3r0fiyIGbinC21FSKeYK5S2VT8ltOD
Dd5ynjexixJwR0VeK4E5iHEQx/0+hxlBVPGSwhc+9K6im6fZ1YiIoYHNREtxr1B3dmT822DMVxaf
iL9sDZVO67OQkR/ZaFyXPNWtLOB1m40Z7E9zh4F4pXJSg4LO1xPHmPi876boUXWbHQhJvWFLmdkS
1lNZ+C7BuyQcrgVw+4ChzKRXzhwY6sgZRFbFhSdC3HkqreaRllAxt74tvWqgiN4EOb3JY5Q+kXz4
C9fx+qx48UtSSToE8w+0rxRuTJPqSDvihLcxkmELu4atn66BozqoT0r0B/6sxbKv7ixvFJpyow9Z
0TpV1NIadvQnNRF4FrM+XC6W9aKlJuevKIw6s6tArxNRjsIS9LAqzKFZCYfS7uF6xAz6u95bthTd
yFUw9HSWbY6pcUY0lXYQRdUvfNXhEG1jndkaHHN+OCV1/ohuHCfGzpcciAjl2sN4DElaBphIvCUL
/ECpUmfJuvphBAXgtbrI3Uiwg3tiJGCf481zuqfwIhFI7p9zCIc2Vj47hn6hDFy+Kf9MYLk4pXyb
U1kka7s8q11jhdebNjMYCt8Vlo5bswGzL/1B6GGNCNrqBZlc1oOJcNAcTinVpi2YumheM9kHqCIX
SAoQtUqjkhopYIBSItw9rM5uyVLX+sYOi39f7R1EVRmL6OMal+91I+bGSyJMGsTsOO2D9i29tSwF
G3o6jIvevq1JtrajQu1P5QeDHyRu9BrJLc6cnbGOwnjgh00U39BCHZCtmiyuXO4M4rg7WLHT1+v0
VVypzuQKwHaz6Q+K9BPZ/X9ASe7fbSSfC8dmYMX6OX/LPtv6fl/RZqm2sjPIOLBGgi0LNaaN8oso
KTB0APssqaaf2zMzhiXQCs9xrjAe7NNpPp2CI+kCDWHah0rYlkz2oL6YqE1MQqRPnquZYtjNQePg
Z5fzSxl5zC+OghwIHyhMheKph5izzoAFu7z1MQQOKcqaik0VQzmZTg6M4nJ8khqZGflV21jDsROD
OBQs8IbWuq98DAhnu81KscorRrrsRmV6etDpKGGzrcGpToWjOBZpifttw9srLuojxXGXh9BPvYI8
Gfuyynx6ahZdAbdGLZgGwJdIf/KSASwBcA1OKWKwExBKUI7Z14ltcHf9I+aT1WHthTKGxzAVVFNO
gD+7e7E9VQHmeyOOJTiGfr/7SBAB2qJgr2cmU4OtiZsbEYKNAlOJXVQuPkkzR/ltW6B+1X9+naDf
NT2dTo6zMf88dRraOSvGvmKjFBqcQ0wNUo+aR9sh/Z7IcWNJ920BZQecMRSBB6Q1wya+mOiYr8l1
muc8PIDAfWHUFFI2YyqEI6k65hhAxZb82+ZfJaS7vQxXQvPMI7G9lmhVLmmxol8OipxzbqD6eX9e
hIuIfgXtXgYTvYclz4Wn+HeuOQXy5MhU4/o9h7HsgoprC8XqVxsHtCEvBOpStSEJQY6g0RsILO2O
nUH391PvRwLpC9WbAGoSzIy1/ZSQCUXzvpEeW7OvFJ243az0Sz+PWTHoGyn3MvJgm+AYk+mvFfB5
66YxBW3K0VxdgfDrP/9+tyaBDbRzE3ccnaERwb0lGnQRLATh4Rq0MYqmzPW1hguZOif8nHvreDeK
BgVNIM5YBcpnJLhO6jeRm7mJ3BKvCEAyQoP0NgJZ1S1n/j1Avllx1dCEpQI9XwU2Tsp2zzsCMwHS
3LKo40a9ex+5HhsQ7vRH0kep3d99hGmcQ4LPr+Itba+KmZp3114650Ue474azYSCXurZm8XizOOM
FJ6UT1+sf81ZcoVd8SI1nF4ozkDmvfouV8VJ9d6BsDLTW+dGvcGdwFKDp+AAuUN7wVA+vKfK++b9
QjN8HTeVix5yW/mh6BXkSySSDzLgxqu7asCI7oTvVAFZ1m/1kc8fEcjCPi6ceTXsjPEI2eJkQLqT
tYgJmSSgmvEBvIfQHw+Zsx2lMHBUFv8tjSv4TDCT7i8TWusS2LrblGSdzMP2ihrrljTs1l69D0uS
Wi3yTE8fguueNC7LX4liPkkyPc2iRVitMGwDnI+2ghx2jgqYWxJSyyLCcVcIOetwTKz+hScjGOFm
6jhtRT9gUJjerGbR/20PfFauTSxYnY92fXAXQ/KNBquZVWRtB5I7tS8S77+wY5qnov9l1qpZjWvj
sNs7/YUoz1/+H213/RI2DJskop53FFLtfBzYeDTI1YxAlVzNE8mKXLFtGE2LwwujQtawkhcRw5WH
7YMYQ6gV0is1lCCK84HaqoWdz3V55Vd9/ldSix0Myj3UQgV3PlrLBRrE1XhI/+LUCHODgnIcc6XJ
gn1c0ctRHgje7reFB3DTq4JXSgfV3nGCGPZHDogcBGCrb/k59ntiol/AgHPwE3+skhWYnADT/Cca
DzNzwAGBQkAW5/Wi6+kArcnOMeszuiIwdKCZ+P2i6Q5O3UktsheCiJT7991svqjBN+N7vaL8idD7
MsGP8B5lSQVFvkV34kkbxyChtD6nmt+ASSyTxX2uzWJO21/fovBdHgSeCRZOhTWPWTSfZgHi7Eso
9F41nO6I8UdHclRrpt79UZKN7lUhKeWBSa/fJuv1mh1b3iYWDCrMkVulGPS4h1tD8t95Jybd23/9
Vlp8MWaH0nymsgcJlbULfvQVZoSs0F15xJ4uMuzrQ1wwtoEP4X+o3rcYwcRmNWSCpDmGWQUvVYpz
5wPC/MK1oJwwttbxscdptZITP5djxWVzAz5kermYriLXBby0xKcahcaXuSw/JFYN4Za4hTn0lYAo
QZzHPv7tsKFFl9XxZSgWI1K9DL7pwincqYa3etksDncy3GHQx1WJoGxqw2U/LT1BH8SCyYHcYcPT
gwY3G6nHAhkukMq4QKH7N4C/mxHcgnPy+1oQHlGkhO5Bh1fN+nVBuSLkrevapSAjt64//uU/A0HU
0dI8+eIAmitqImNP9cWdsfERyhU3HySDKkISiZV+5ANTrq0v3r+ORhT+b2S5Toe9U9ePLdODR74Z
awm/JQ1efGxHm4gLo0vP0oWqGLon/aXG+TAvmcmjgOr5xMyEpG2qgNFdhbOZ+I5uiP1vPdF826ye
bVHyY9vIxRFJIzXJ9dvVBLaLLyoLy53pEhVSsPF3ti3uCIsEpg/FsMcrdROlD1azQvNDYMnOAyQs
IkDAFrZ/hc1Q4D2TdXY2l68HmxupPzb1yOkkYJCj4v880uGLKvxX6gwkvE3KWXRmYfXSSPP0jI8e
cwdB1n/hdYc/Way9ajX0M0be46vj3SWl06jP5+0c0RDQSRl1xPbDjaJlVj+TlM2tq8PJrnKz5FQV
5WYMhoS07J1PLKoSPOZxtJZGS9KVT5FKuNIfIK8RyfJFJyVArQPvJqKHUU9PsdM0QEGWJQ7a5ciR
uigq/YrTf2tBh8edKMMmzg4g9Pf0IZKz97Btb+1jKNBN/6cMpthPL3Fc00Zq7TfpVwx0u1uzL07T
X04nSPRrGLlfl0Wn8KTnpGjLhsQ0s47x/jY7QCRmjyFmB0AXyxa1CNBLZHFR3kgCly4KWLhtJBXb
lmh9lwOfsowjIrin7Z0Siu3Ezq+/7qmjqL123te154vUVjOgsVtJXgE2iNLMpK/z7l7iTOd9T26w
NVT8MuS4Bfz2PwJpP/nk6+tNuv+YPWY5n27cYMNDuy/jwZkqrn8vkKnrB35to+G6fMx7mmbPeati
eSTpJ4YIfYjg6GGJW+Xw7xmUZojcR0eutzHBLW0pU+kjJ/UdcYHoqRu1F/CfbboAZD/mlD3zlVlz
1+DfJQY4SyW1BT8VPZ76kV72qFgQDi+9fz5PBWi1SwwipwQCIAGmOGMANmRZwmeMZsHp9F6bf7X4
LtD4WcfiKMEoHGu0t3dAdYppIsL3TVzsQgrEJqJl19zR5+kBYxu4q3MYS6hlpu86omqvNn1jFZyD
QmYDb9ZlrKADCCcFrfQteDDEiZid0r3Pq7DCduBGHhCAaXnRRVghAfD0XLbhJPyO7j5kxRt6UtDq
WWjNVX5RwEruU/RdlanSYU3lToJqaPBR0aBqxCVnHN0nQK5WVRb5zUtR0XtJJYgZVUyHBhJgZcB/
JQvTuqe0HYD8iUQ0O620kamG9KoAFFaXy3kzvbmiyp0G/K3rqufSGlLtUxB4uFi9a6wF/uvYmXFI
dr1mTgX7zR0nchOiRmlv8N6kpbBJJDY/wG0cHLAmw2hpDniTEerL3JKZ+UfT6s6sfD97rgVjLhEf
xGs8YxcDcS7YeqzrYOIGiQZjYVz2eUxHtLLxtRDP6QEHzuP2Q21Xj+pgkUHE9uws8w7/MGUkF0o3
ajb8Hq7Ojggx+6SBkxAPXkOKX3IfJ1Gvzm457J4jiIKfraSNxN6itSC/seOREBN09je/CW1q9ga0
pd4oG0Rd0Cb3aCtPyh65VXi98mW/jzEA6VjGmEIxDFFP+PIg+Q2fWptsS8ov8kICnVcEbT/khKJ+
Q50lkkCkuuYxSaHh7XV7RPIaZVYqA2xO3gBm6+m072Yi8ptHix9AodDJvuq0rnen5WiyX6CGjuBe
xrd+XPrYYPxqXI0i9/8qiYYpzhtYngSQ57dqyhEa/+41qeKGBCwybLSa07/m/z9Rj06RAV8i/vrf
+x59UydDNidNe0KdGccvIHN6lde6PdG83+DTQ6LYwuj4AW/fCdgGs438e3qug+b8C6G0AZ3SN3oS
La/q4veyR5FjhzTXg1Ub0Ju9AqeeRBtN9MCGdBb57PqEnmRwAqoWVgRWinwZVMSWqZsIEvu7asie
pi+IQofa7bCmcJtCMnLadM+t02CGuRFMb4jHcbZRw2HN2wM13NimUhQfEYxAjNQ48uQGWJcQiYnz
i3U4Bvp97YPl7a5zoKZSI2UjogeYSPDUyHR+31N4ibRTHO9AqKP2vhuCWaYhbjdryxoMzd18PZCQ
JmuyVf8RhivNWJprGvMCDx09glfDaa5AerLTaluDZ7eOydexsTNrzgp8/QsKIBrCPCdaC+DjC4vw
8n7JXLtGGf/hpYvCX41TDp0B5O/Qa0pFoaCAyIdMjf73eCcFSmJ68QqCV3w5J8UR4JpgJlHjHBQS
11mtoPiE7sFkdouOJd3brFLXak8WSQuJJdleaUP7OT4DJe0R6IuJJ3VOnBl/fmyTlUxkoKpKHN+R
VkkfP/0K1jSqDm8hjA7/nChpGNBweOIldYJqKhLiomYSih+kKWcRZcWJ1ONRWY6CQp5iSfhJoyAa
4Nb7uIugIAb4gCpeZ9W1hww5nC71hTCxabLYRZjaWUhK5QikikbYKJCbQ9VuCYS6fIK4P3LcZO+A
iKGY/UpzfODdCRP4xRLTrx8dgbLu117OS28RQEvlICuLZg2EumS/hmRVFHQ4a6EkH/8O1pzpAi5c
QtE2Q6WZl5gZRB4WEdLy6VbCKb+I2YywzGIqMTP7EL4ydBd1LsXXbxfOJHEqYTrp3elxM+1tHRMo
7jRmGybrdYVuDrvpjZX8FIxKblQgE0w/v6413Zh3V6HSaXx43g8kL2twgx6jr5e2W0Kkh0Y5ZY2/
ylChGTBVmrU6e2n+rVdNY+b+Bw0pn0MeAgvy5ZcsToAyINhJtkojPWpr/ErHA/XzLISYY7vVWIoe
6jT9SQh5C6Elp3pzWHzDd5CxIDhrtzaWC8MUWo1Q8MWBObZ80qFgwx8cOrOlYbTuCyIwA+opLj0J
wMxOs5aTXn4KDe4qz6NDvlAjNr9pgGv9MPip60FQwwYHom2Nl/OHrav2SLtFOpqLxGsuCxswjXj7
FhXLu7fo083JDXmy3gUwGmTnnUYMGwoNQAcBUtp64Ww0vo7zCXId2rPwBhdbSxNaPa4tDSo+6HxJ
hvOxwD/OscFqZF8veC2otT5Xo2JKypafnfAwNeUQE04/MJoyKKPSMJ59qzqof1/SqaFNGXEZOBk/
1uT/OrLtugZqu22TvTBvjLUXJuY4G/KGYRcxtOuhPel7P+l35UIOwwBRVm9UTg1Ychiqm6RWPl5G
RUDJYLmmZudPSqCmg/EHoUEW+Cl+QDh5/QryiPTSTc8Qtocl2+gv+y7xKRhV1k9lTl0MIb6qO9ij
CIChe7yJiAALgUqheO/gh48CKyTc+2+jjYXaQWK3q0OR9mhoAPZqD/ZSoFNg+P/OVNqNgFWQAPrT
LQkfO/B1PoGsSENOJV6yDLAu1sutj01MsLHgGYHQz9Eynsn6efOjcZkCxpO2CqbN+FRXic3Jcat3
cD6mVGHIctDuyEsRRgqAg9reaRjU2gWb04RYUMszOLkfUIEmmES+MaMvS0mrw968vbju8DE7pBS5
dKdW9Md7/3zQFjUjHib2bZ5KcYkWU2pUyJ7kFIS9Ow4ssfuid3EIF5ySYJvkWs/mWBnxiVgYODk2
zjrHKfYAXoaoSFD6T3RDeX4WKHIBwFOpg1VBILco6VkNGyBQ+th8ABf38DPab0BLxHLM0Ti8P147
iVSvf14iPPxgkkNYRWYOOrM+peA1boQofxPPQslI92RXRZSaS5s5dkUvFYPZW13QINrwEJqDxV32
8X26alCmTG+bsDAFSpFZ47Deve2RN4BBSzF7sB5ct453PKSbW8vDw0OAnQLSdsun0EjEkmfBZE9J
/SSoFWQOZMahuoaOKIBSm7tMO5RLH+Y6nncZQ8evizlyU1EX4IWL8y43fALtRR9MSkPdfzxiG/rS
xMH8L9ByBzC+r2jFnTJvlW/+O4+1lz8nRxMykWfd8BhJO7ItzPVExnBBaIOv+lMq84qBGaIOgrkT
CdgRgAaX6GgqtgEeGCA9bvk8uTbHksSMOoMsN+b3mc8l5/sgcCJG4BZP9luupRXXGWRKOPp0Mk2/
9QQAMCaFv0SLotv66syOuGAl5fXHw2KMMK3gNdgprRZZPT4r2kdrOQKAO6SjLekD1BEQKet78I+C
J77TPUr88H8n0JxZlv6OnwvmaIaCOVDKvMCHpz0Wmd1piv4cM2vwXsYQqBIywYlxte1GHXztgtk3
Xq6LY60KWdMWP47QG3GikTz8+jcB33Eo9ynYsf31qQ3csUqyE0lem2Kk6qnxSOucAM9GYRAeB0CO
8hGEwcCgSO2jo8NBZXhCzQhPQpDigko+lkb4tCYzeLm3qARvHIDetR+nTPx2ILGX4YDBiD6GXDuk
BTn2O0WuX20QqJ3i2V205XgjPLgfERn3UkBTA5X8/WX0YhXcO//bpkU5cWqcnG6RgCxLl6SimZ+F
Cpl4jnivBePInz2KLs2qjVnTrMfOTzSpRvGKVPFtEjh8eIzTUS3qLJPd8U8JQFfNjc4Qu44164JV
GxNEeErQCye/vWqfof81KnqhTPENGvriV0ssR4Pak/xzCb6r99L1rTLPJ1dHVAJVDiHzno7k7vxY
FzxY0M0+GkLDwLUpgC828tPK5XbWnIztwUJwCUazGDwPvliTkSy5C5rAUqssKr901TgHXWmC65vr
w+0yc+YJd2PAU8ySDWZWtEIDxp74rhx4CvrVeSJsfplykC0YDa4suVcAzheNTb9a9QWBdjrAEhOk
HWRAjdtq5Pr47FNUkVlDZKWzAWl4gR72JUo6CoBV8JhvT3U16vU0aBEPH4KcD8veNGWBvKuCKdQy
XElvXsuhZXknCdoMWOBPEUv5+UuK2XETTciCF+m66HcGstAjyPQYYt3ju4y4ZIwp2VX0J4ElFtLA
EopRIID67RQGtoP4cn/PRaQaIRfBJz4bMUuG0r7VTM7919TnqCEg2j+dPY1ryum54ZvXJwx92IDx
O2XK751VIWR6bK2GOA5vs7Ryj/Pm1FcMySJW5yorVt1s61qut7+baP4dqdYHsyPM4VblWILxmSk7
AvceaSDaMt9pToR1oSBo6Qm3Whp+KRPINvFXcOItHUgJa/tZvQAI57V/MNFsdeqjU2zjuGAreTKH
FQZzhZx2tdpxlHT+nuhURKR3HTRgkCPNmHyErkkad2xRF9mRHMq0UNsY32m60dsPNJjoHIGv12sp
MT+T6QwdvUifP7VLIzUmngCBfuQfHzl7Tl/JSmoWLk9Hk8BR92WXHTiatje63emfJXHUj/LwjlJy
VnllyHNsQOTJufu9rZbx0S3JGXS2puSm14MZLxZoQr8MTgfIC8KtVqz4zB20AKMnefowuewxXJ/Q
WglXzVDcUoAdz4SbKeGsEDeDeQiAD+hPn/bUYplYhnHsPWhOKoABCtqNmScT7OhxO3p9AhIfTbz2
YB8Ys7ohhTJqM0/kP/877SkDMEamtwaZOp5tgClUcKWjilaRhYe5iVNkHLO33t+MAz+d013mt53k
tO6M4G9sh+WHZ0Te9T+75LMUjavRfPQScDZULOpkVLSQtz/XGDD8+O+HUbDaaSQSR4rLe4D8BN+F
Nb/1A9gOFA9dA/sRZ2XgKdITtc4Br6jQkteAv3ACvjl+fZoJBQ8EAj7bcL7mFOwkmuusbVnvxD72
RQbFSDWzEloiOKTjzzq5gJ4JX3eSMChOP42lZckdcLK4gAHiopIxWJohHicff/I1q0RuWq3yR35d
k3SSmUHXr+WP0WhnUo2gas9GTJ3n/KfUyIOiFwbXc2Y/suMBhMwq19L49cKuk7eKWrWS3ndsr5J/
xGbc2nSKzsDbYlOZYWWaAWEoXR6Zox68WYnOxBMtzDJpTVynAgYs3Od2HF0iToOV/tS89Pxdq/1r
MAOFq5NUaZJUwNKmw7lB1DsKZ30x83b1OO84aGpD/jpXmTxsD/XPShnlTIz5splWNPfW4ZpX+JlV
GfaM2k29/8GyIh8ob5rfzriGaVMreQalD2cs2S62kPiTC8HmYqJKyAwhz35sq0LURZQMP9AKNGdn
a1DzCyoa0ejGdNT5T8pw/h3eSieCA7SJv4ELp2um4cUvFbFFaYktPyY65CKDE6R+l8QdCTWw3JLg
sT8QptaUEahyeL0W66JHtpUqnHP39Bzj0JGgYpEcmugjeTsw737UZ7OgZ0iaXY70IH1ZIYVCT+WF
ZklA3x+C8cp3kWC3bydob6At+oTEeMrvG58OK/3ZaypkUckglXin0WMeAn0wLNyk5lgb/oYULCPn
DLlznpfrSpjzkvOB9JZURahR1zeM0Qy2Q9gR8f861LzfViBaemW476qd7uE/lb23Kw5dTM7tQgNd
duF1nRAtT6hm53VBzr798pnGh6GOT90nN2YhaeyWVfPueX/xImNMW0NTksliWW3E+7omFI/dgasj
J0yVZdOS0F5U3/h4RCPuj0v8J07jQclDeqmUUFUMVEdeZ5nbRzYLooLgYZ/4o0AoXm4zPFvv4/V4
TDOPPs5tcW/ARwbr5uESPP6U0qvg2h6s9YV6TjOY3b8AZNuVS38gx+cnoYKrmG36b34s7EQorbNr
Rd4a0vFy/axPg3Gr600t7G/EqcB0ZR1Smq98AzUkLNpzm73AamTxildz4wOmeyDNEeRZ6E59k/rK
wF3V0eIEtIecKXivB1KrnezRHTFZr6aePH4mbdWxPxXfqVaq1LfveCE3vSqDjY3qBWsMCjYSwsJU
a0hsMYG5jNuBToSILl0OaeS7ruEbqcy3AXwDO09IpGG0gCrnehH9J6vdNQ3hAqt8bdw9TOLi1WUM
iG7JV4FpzNx0RskhH6jtBY1Xh6aIWHliZqrMbIyzEDBxX0Uq8Cp3UgasQ7LycpNBQ9lw+kxkDsWy
5RABuArFLmUlwToAnshRt5GTSJUrzpwpe+/L4aHIuPFIexKXlIqcw3wCTngg/zCMm3731AGUaTua
vOrQYz+2Yk6yqjeMeRks02blQYDvTDE8KaWlGcCjrKkG6yw2NQPeZF8seIltYZ6m2pnGKI62w8I4
FWZ5oGlvcyrpMqJSI7jx8PjRjz30hSeAFDcPw5Ut/rzweYxK6tYLYKDbYTJgMVKpU7EvVINv+9RA
MBYdPJjTs9K316tXAXrRPhgmSZbGdm7Xo+IwRvKKmOrP0/S9nwxvDwc5uPEhjCodIqrUax53Go22
AyYPTaPm8vDTEJTdUNLcHEIH4VS/PDqYyMkarjSVkDSYAgGAiYgp6iWlqMNuRFrrxsZCbuQtUbV5
G8sgBSdx14GLIX0gumDhoAolZ39h+EHAKAInRSbfDDoBu/jTODWkeZ+XIFdqr7tFa7sXsuQg8WbT
ebDKpzD23LAhnnnM8YbD8ries7TAKCmawyzyaZF+MHOAiJRgoVjL+Ep3u2k1AvsxIIxD/HTRFokE
lVpMB3Jw1gpuziZQRoxxXeP4Qvc99gfr1gRdlJrcXd9+elphA345M4TCsIT7uZeXYYw88GImgMgy
e81ksCkAJuIFp+IPD9Ralke8TD9RVfT14NXX4HCZ7r0KhPnmzcZqdfwZy7oN3ZnyUwci1Stm3Bq7
WMqmJ0NmvjxDIarvO30JX5nlhG8dm6n4kGL2SlbavodktjNmbgZgtsi9vqMHXtg3beWINqSACPet
EEqm3ZqEwcP+YLM9Sxzjfztq56cCJS+taSrKnyNnO43xxFuqCh0WQswjPXNXIbgWpXMsZg8ajDIx
pK+9xGE3o2gYi1ZIX7vcUwTGviXRvAOUc6w1POK1rVX4COA3xoW2FTUnTyxUpGbHwei9LD1GhCuR
zzPdawVL/MFTp+Ng1B3E8pdw4NpHz1z0QkFj8yMHY58WuIi4jtHcmoeHP36u1ln/ybYVp8eMNkJZ
lsdI8VqMl3EV1hwE6iFBzX1mCC/S8PtYNooERtrD+QD+4kpN83b+cnhhZkbGEk+RPrRKufDMpjuZ
8zDlIszAo+FPhWStDptT49T3wFSGnaTu5RFJXn9FJyXjORkNrbfuMHjQG+toUqq4KcHNIgIMYhdL
DhsPKDDhub7FHA3o8+1se9AXCR3WmC9if9HQUx2t37ZK+LjVc0XfsijQLdEmj/VDWD0gAiUbyWqW
3ey6Ue9IrVHW4AEBt6OSIMpX7GxG1FWafRR4wxVoh7uMsi3nNECCz65LqL4DyIwdojxOplxBM0Fd
zwrB/NYFhN/8sH/9vDrxWmxK+qsl9mkoWulfrFp3TsH/0TWGaP5cC7xnYNdP+9+BDEXy+5mskMCO
m+sHTXb9KGZDcIsTphzOZMSfF3Mr52mBFWAL5MT47/MbcIKiCyiNTU5rmRIQsM8idh3ShVaqPly0
SokyTaLxBFodaFnZWMAyY9NaxpoTB/59MUsOKTT0cd4xRVPMUwmUuDsrMxDG6UKRXhkcPc/XPJE1
MZmx4VtEEtK+FTx4GglQxWHTERG328Q1BJoKwsmu7uG8ie2CCEJ8FrHyHcLfKxEZ7xm0RKo67dYB
1O5y3zp3W1A0ZGbyAcwIZPJlcsFlL8VnJBUaklOWl/r34FV2SSgqeK4GcKZpTVe5SFkV3tVdWa5g
KdJwol0Dr8SjmvhpcPzeXyAxYBRlYa1/q8y/zj+JbkhkdoTff8YFAaLGunSRJJ6VLKBoE5PZrdsQ
VSM00QM0r/QR8snZrkK4rNQcPk9jTs7RSgFkJdOypM/NJXsWwH13HvKF8JXSEHPaGob7KaxDzLPg
eaW2GKiKuaXkQaPhhp96xtWXHta4x3s99PYSUL2BTWxDu2VNtByWmPLHC7/DGnytp6o65TPthnOy
JvNrHLOaC68m9xgbriPw57K/Dzp6368WkArYqWzazWVo4DYmx/8RcWid4mFCyv+SVYXgPmxFUN16
IT9Yx91D8Vxvg01TvXay/zcZGqzPm4ViT2al5WvCfNd4XzLz+/8rud1w+1DaDAqriAqlKXPQiom1
ifOjeFZ8FZb2orMvCHftrVp2CtBNiwKFMK1Hz52e+6LrAmtxY9UoZU6RJh/svJ8GCIiiPLM8Umzt
hFGRGq3PlwQUpH/TPnAFX8zTSssQaqvwhkO+avDiibEDDXfvhEmCwMRvzjQOeMPdpBrBl+cx3RgD
Zu85gnpatby54neEc8D85eocKLG6qByNJgqvNpf/lqSMA+mti0flMRPDIPNiA9Y5aHfRhdv+l7tp
QHjuM1tvvifdH627lDzHyChr/RsW+8heFYIVbjmMjRJG1ZhCfjFlHIOGK9Or1+5EYC6iKaHciMNq
dSRIDrQjvzeJnkt9wHzGc7aWdHzuUES1pofbowM9tYWMWrVxqHQjPq++nYBBdW8kXE/S/Ewgd9ML
FgwWaQa7M2RdCAUaa5+Uyc/rC9/DIEyP1+u1UKuR0XIg96rbdIFJs2P1bHq9C4OdjxqTzBFjFn6I
CtNGZ99mEhfjEXuOamf00/PdYn7Soruq0VDyO1vo6OI+6FGIv8p8OXeMkofnyq4EThtEsIphOVAs
dNTGsqgp4BFS/S7gAnsdtabsQl5AWd6hHMAWJsVFoA46hiNYeO9RQbJLkKZX1Awtjf4+BfDIPvtD
7w7maddpss28pXtzNwJwsRJ2HNSfKBuV7qBighdOaO981gssu2/9m2s6nXDgdgQ0p1oAboWzxxFq
pY9XPHHFBXnXuEwlJS+Z3msu/y1gJAoSHtD3p5fCnd6dnBqSETTmd7SdyYCEK37l+7/A+8bi41Nq
kIeTGfdlKZGKUe72ybFF/3xY5vdk5evKSV/C4yfXfRQfgUwTjhehOUCrXAAJqEZb5AGrtX6zTHU6
WtOXNEKkTh+thD8sCF+nl4qXyusdav/hlVYDDb6GuE7v9dLzTMI0Jnde72o3yi7n7CfuqdWAyS6L
y0tT6prXMqAuNrovBM5nNVGeNlohxe/loy+jX5TPCalXVYF5I+gFpcMI67lWPVWGl7VMOuW+EYvr
Mx1/XkjlMM/YTcAiG1DVZB8ZurFDdDRc7KDKJU4NgCn4oQA072Xi+a+lKS8XIJa5zkV6RhTcEpQy
ErkfLlFBxgEMYbQDSPs21EKWz580P/WnzoVEOsUGEHLKj2K+NJJeuiTK8vpqfuKxh3nkyzqsbZoX
1gLR6nm8riOmvRyoItdKoVOJIdbUfv2f1Qn6goUxccTyIywkpL/AHRT5XRlhshlUd8idhEyBJqzq
5mEgTbqnGiofX68iwBrtw0kaqXHR47dTPst4JAVYUq5WZo1jEDG94AXuSCBeY+yn1f8UO8UE+kEw
5BtDuvFwKSBQWBd0CRuaBtUoADHWrEb0xe1g+uQpwhd1ue3komCnFhRuMPaeaYiYBW7Dv45JtZlc
CvNayYDVyglAy3ZHNncWiZbI5Fwp2R4OtqBIK5nPHeOFcjm+0W3s1rCUvDnmqwy3JRJBqT/ik3or
UMmSqn2fbr7c6jr2AFxCnQQkj4HtZPiv66j7nVQavzH1Uj+iI+3iGbNFYMgvzS9CtoFnso9CLdK9
N14JrtQVhdm02aPMsXy9L9c1a+dvpJdzGsz3k6oJkjhX0fQsv+xx3FRcJYEXRVH8OalT/uwxRARX
mH/mG/ibRW/f/YdELLNlMG9AOgH2iXtBCmGm9riY8HyBAIqUotKfi/2OAe0sygTWI46pHgCdfkwq
bMgSiJXEzHmo7N9fsFSKMygJNR/XNGXE9/cEbfE62TnNacvceIHbnXMEn1L5pphg88iNfuwHE4bY
gZhn7xG5FpEPwfHeFnB5TKoFsJnJOWvPqmrKShB2hcLmw5/doDbF3D6PH3+47qZba4+WNQYA4urQ
azGdV+gioMa7o/J9rUxVdASHOWOq9wnrIRuHbLuyMsakQlI2O0qnTmVeUN2wAqCtgaweuN4ucSN8
TJMfIgLQkcr9a1xielnwlngITF0ucbr7WnOPanWe13/jLGM4pf8a4zJsjNXPIKBMbAIw11TDPdsQ
Knx1KsKRaW69uEPJzvJTzQR4rn7XtG11owHNLrNL2mEhEuUCt4DmP21FEzgdZAFG/luFoINhczca
SRZhbpth/dPgKa87AzvmqikCUO6fn17ZGhcqZxoTBUCvtSnglhjObn/3KDuDhSny9VDZJO0dihkr
nmI3lF8UtMcOjq2ffWX6JTrUfx3kbMYgkh0YGOR7tWP8V7V1SmZp2LMGeMTxhPobQ1rqEKozSRUz
0jFydWnJC5BwimrsxbUVc65GVAKfxSHpVSB+pSNJxOLWB8mJlxhS9ZWFmVB+3+nzWBm1XxN3UQiE
d1p9Csa4FeByqm3us3GLv44YEu5I0Xe5QNtEp6trUJcV3Y2a7MPIGUDr5bdFuOGwj1q9b4wkRWmi
YeJA7CCIcnzYj211+yyoXoSK2wugYuyPNdpHKLuGgBJN744DD3pCBuFG1JWUN7nCDPzHRL/TaoE0
5g10/yY7wAK+XUFW70/bZoPO2Dfm4AweiEq2rqgefhXC6Dy1b439zuMV3KlD70+aEvo3hzWir6PW
9cZqiNHgbH2iUjZARuxcF69hhgi4CeaRkAkjJL/ni2A0TPl+JIu0y9VSAlTdzuzRCX339VST/bzU
1L0FLWNfhqfVv+f5yZ8VqeEDVaehYfiIno+h+7LneaV9tLBjsssg5xZoYCLObc+mfN76GJ6fY0zs
VUtIoOZJaEC4pZcxrU4BqRGkf35Q+FsnMbtQREEkM4FUWcu2DqfwhKQ/UZAgVm/28qP/CJsXExv6
RK+qNS+EBAE5tLDSssf8mUJfX3UWJXhSAQVl1GFsZWow9GgcQDIo6kgguJrR8Wdym3jDjan574fO
w/ULQ1Ag/sMEkmIp/vB/pD1zsCaTm7Zq2giqaB23vjPoH45RMH3triDrRZHGxpoDlbstnuHCAqg9
diijPTRSq23U/QfQ3ySZ59Q3YKwW3N7DfTKrU2XV5ntAQUomk7qxlc7RKTAmO6mgquSpz4i4pf8a
fh+DpaRdAOozerLYnrHNo6U4Up8j7n4k1No0a58+xrFK5XN27XAw6ITrn4lqn5VzG2fa5LyKhcNI
EHQcgPABpPf0KwRhzcmCz+ZpqNumzEYZBmGwpn9yrc9fbTZhsq5VE3M8d9Gc7YrYh0biMJMWPbVI
rp0/Dt87lLoT5oY9LpngNB0f6h/Lc5Lm410cYyPOYB5py4iTelK53RyO46HiMelYfuZXn/G6CEmg
XAghVNxNJuZuKkDKFh+fzr8yxc0hiY4M4X4PKeHfVWiwZyBOcQXfPglnHLuL1QX4N4gg7fdAPYWK
ENPm6PyEQvcbSi6RcXSX2wV8q2hds9MGBQfCqHBJD5LIXL9NOI/Nlh+enEcvTj3aYll78FiYuTDT
MX+a93er2mcWAt6o8EkkZJ0QBcdvKCibU2wA5u2mI+dkQMzG7Qvph6vNOn989iZG8OmJ/8zjbzLr
gFeVIK7KNnDV930lbIKcicd+6nxe86F335CfOTbvujnmHG/ZF6ZGje8zuC56dTCtZgwdDNIsBOoQ
HEGT722Sig2aRVL6LlOabwh/ImXhCagLOrn+PRFV6fyS/ch5yo5lvyGZfDs64CfdE8nRjwytmtnG
watxk+B5qO+wkqS3mC5DTy8aIbBjMVZsSO50b4CYNSQZAsSycS7UGH2z/QcanmJOA+I8KtiDrQ6o
nLbmDI/qb8PimY3qWxfMhXMtZBOaFUialuV1D1kqnlR2acqe3iCUip2NXUVFJJWcfBwnkT5v4N6H
ObHx98qhTeBC5TNbzPrWf/bVv+Lzpu4PKhOcw3bxmq1XecLCo9tsYLYIISpQlM5DaT7sZd7IpuD2
KJB+Q2znTOWDSL56Gr/Pxf2G+TZ2hv3ekqqf9Aby9+xU2AVaKH3xn6ztURUtWHO/KL3q3HLk1eb/
3b3XAVK9xDjr6PUHp0VmTZm3WzCSw5J2mSmyN2uHjBLttSTbHtPTxH8Lg6vYNmyQ05GczKhejWHF
Rfyg2fD4xwNqGw1Cti+/YCvlKahl6fNgSloGAgS56lHXnGqjtpAvXoRuvQcmC5dAtkP9jX7vT+86
trabWSi/P5m2FruyDMaamKopm1L94RWPNW1J3UFcux8kJb245xe9as+MFF/vaUQYW7n5FCPekmFv
KUiYJjL7KkHJtBEnd6GTTG0V1YVLC0glGL10i/OEKiMMPN7Pef8lIMH/p1cSJT9TwSyTBlW4n9bb
/6gzZEp7ExKSgaMgxjDWkY4d3iHwv+R/kyVWM+qMRfWAA0kTe8BaTKL6Cf9YHMIGjw0pDtNFphQr
92uGHrvTlqsH1c4mPy83oqxfWfkdleFP5JHbJZcNHcOKTa5Xp0MNCTHf+osyvOoDqq8PjgQkwqjF
BSTp1CmzurIgxv7iDy6tOHfHPL93UcBdDwEpxnxLHtIRlfrWawYU3IFiLM9rhrhjxj6EkuFu0c4Q
iascSOQr4JFV/KahowAioRXAeF2hl2VsHh16iPM5VRCEZRx/3wR09xqv+sqAqYmaviOnY5BFnEAS
zVem3FuatlqdDTYwkQA8Ct/4FDY4L2emWtG4Y+oDEtPiFOu63s/0mTywkdMJvfrSosXaEbJ7KB1+
JcBt/+uyXpfq7rcUJ0oWqOTpbNT6wyJQ81+0k21eJrgnxDZIcZv2MPnmfe37AmtreHivdQjPKjsS
FravWIx7wwqaCWSArwWzQo3QgDllb8Tf7PipI4dhf4belS7dHs6hSyl9KomyWfFezzXg9zxuw7Xn
wog1CJINRPfZE+fZDkz0ra9htzf+TrDAwscPdlQrwLJyn7Nv7I2GyScBJqoaIHqHWwD/ZBk8k79R
Fw1uTZzZOQ0vpKuJHGmIRYlB/yHa6Vvc3/p8FiiScFVCLC4glox02WONCDPfrbPsHbTh6ZjJcaY5
ZfzLweksTBTzy6XO2qnCUjnFry4CiuAhJF9Hi9GCY1HhaId9sFD+fGwhfy2s8EJ3TTvT2VE+jsAY
npACrpVnDGrbnsZiUEVvnG4XeAvbiE+X7eP4byjUSLDuBWOamzXdkKqYX5CGu/61+QXG0h+1H7HK
pbOl9fLGfwCu4I8UhxRrDMPdB9F82GaUJ0H8kwfxC3/Je0ZpI8hyb9XZ9kKRKnoGeOcWX8IgV1A9
CXdU64yZtmpCdfDYEqQjKUSzYDlVhoRu1cmXISakdakzt14Dk2RIUWHlsC5lhFjHTlO/4vkFYizA
EHeoTnoK5mh3XPbsqz2FmGyNsoKisrXj+KNWnoyZ+2Mc9HZdN9z5tHVJMDwStgLmgjHZKmDz6J3X
cl7PhyVIMfgVawyyaOsaJKCGAgpeEk23Jtmp0DEjffwtp0xUC/Agvj9NjI724YuLithl4fXwO60v
Hgut0pu2HaxeJMGoeWImYi2veOqdS73gIhtxBM9j884694D1ATlQ+Jf/tDrMWM36kp2fX+cyT60z
JyNWLvnVJ0WC/VEWb2bFdrpeqh7CQLmf7wGG+dY3BfOg68m1XmsYsN/WFKSUFIHlmvAO3J/lHDXz
JvBSnBXRV5ri0+Ijc6Afyjan6gp4agT8UhAPiCU8nxEbDD+eV2P1ALBoRw8/fEmVQZMjwlOm06y+
Rf84Y0iP//ZjXQtZ+olsyE24yujY/LydybNyDOBCgT/bAb7NJfFjdke+oFTQUOkkWIU7iYtBB0WE
1S7sHQfOnDj/ZyO9M9UTtwmLhUUGZmZ+0XDzhuHtcX+FIwhWrpylAbBItLZKBMb8fcpd7ueFM4xc
zoAwJ+hS17nua699AAI83Yai189FsZwjU94WR9x0rTeFEJkSU1TS1r2kpkJ3DqWzxZ88G0GTYylg
hDGOqxQyyFZfeBq6RwZnaIX7raRAgFWi1XNDvY25CGUGTubhkX3BU1fB5pfGEy3bRw5VKiZM79Sj
VfFJYzGGWPkzE5qnM8+zs8zGkY5WQ5Wz4SLNJ/N9Zy1eCP7asUkW/Omvw/zddcPlGR3PJswIPrhU
Vb/cwXAcGuHNobE7HVXUoXk+xkvtGDlOU3mWr1LUmAc+UeIzkwPHCeW058/TQYRtaWcLIWSHspaH
OUXW+502PXwy/aI7N7rA42ZbhSQTbA9PAZYuRWQdBYCEUtTqOVorUCKgXG6NTw2/McmLRP/kp4mN
N/YgTQiiFHJPFfWNcm5fX5DfedQ1o84im7P8b32xldehBcAE44CyW4Vl6Fgym3gbZBJ9DLKzlcR1
oiZgBrQygnBm7X/bAvrvy6z1slPWagM57J5dy2LX436ZW4sRUu23oH5agH5iLoRdju5HdCSZoJhd
aCdyAbWBjEOqesLTn81PkeYd+PPuBlW4caAgUCY3GjJjdFhyMT7mRTkyw3RLL70Wtb0b8lme2Urd
BJRN1b4L41tMN538+5sArgqtwpASxfhjonsH4gX00RMy2Gdva/Ygta1olWnzy4pm8IL7WhCBIy/g
liW34TtXOUXHWLRbqJlOW0EHw9TPhwOFpQUFlTgWl5gEpPA52ah8W7nA4ECOoX7brbSp7OBxWyig
s87a04f7kHcMAIWkc5QTWTLx0iygcdsobGsDeg/Z9ys/2RF0eUi7HOiRnh8AtfWSNiZhy5kB0Hnt
FiEBHtBj50Sx8XhQkb0xdNjAyoi8HvptcJwa7q5nlgv1Qd/K+TAifUf/Y0UXnmuS2gU/j4Nui0ZB
HvFvkpr8Tydsq4/YmCxd4h16kLDKx4Gho3he5PVH3bXY4woovH73FAY+hilZrsq4LIGPDfg6dlOs
6hsxMlzAX1Du8sNGRQFzRGRn9GASTm+s6yD7yUaNL2OilHDJ1PgVCeQzw6rvbi+bxMvJcTWjPP4d
0Boxm2XnlXQgR98R3SGVNzTzWh6WI7yLzXHg7GtH4Eii6hsS++rcGjujdmwnjjVVrmOIA3QQGuty
9GryISoawmGqZow6DthLzpagEbQ//IQc8G6FV8vInY/LuyWe+7PSKJxNlZC7MiwEmwKDhasPicwK
f/DX4mTuN2kb+ZGwyTtvuDoEok4+lggzvmtVADUjmtIv+7Vpg7W7uEEIcaVWuZEwpZ075twkChUC
HbpWkC2UIfN6tHE+Nw6cVN3iJphs2ZR9Nrr8/gnkUH7dQpqQOFXY3JxIFYtSk68czpa+6IuKuQqu
1ATAvhCwWkGjVROUNACB/eyA4J92wBZDBTVSLl55b9rqBzoMzewuVThQdNNqP2Bb2Ut6XOV5i3dZ
ttMmEoeEJCkKk1Dt/sXFAGibE/zBemj0tIlCecX2PlwC+j1C/p6TgzizgtIHbXDJ1IQYgk22QDVt
WOGOma4ySYabHuXOdzck5tep6nVGXsysDqR+B+xVQrVRAMFfMHWGPo2ECQYmR8Er4USLhGGrXGlC
ggjW0O3u5lmwh6CJhFEcZuXRdY70JC3sg1X7/D2XKgIXopSdNhRB8NqbR5Agz2GpkzNxBbZ5k/rY
pDjljFfMXsLNnWX2it6djcmRcZ+SOAuZdUIaIpRoGb5LUwEu0aXUQwT4OK+30LB7uA6SmA2wBOSN
QRdhTRpwoMw4yVnTvguARJS/1rqUubh8+i0R2KP8BjZ8CqYzud2Oi5xcfFEMMssb1CTfPhnZgHXU
RTHnWiDrZ1R7byDFLjdWOIPpOdpSBmohNCKs3rj1KU94v9fqe4CsALLOVw6Mppmum3pB1tiUCf4q
k+sZ965xL4VhaiuuNrHEps2D1V4S/W87q7F5ixLWCWQ7J3jQzLNACsTuczq7I5S05Et29Kss4YqC
0f23kI5IaTTvJD+yQOPHm/OMs9vaeuh47P3B00PFRP/AM+pOhHjU0Wx8e6+RBtxbz9kuUGrQjDRr
XrLTyGhtP2BXt1tXaDZLjXiS9mLb3VbS9juTcR9rzBAH15cY9updmbknV0J8CA7Cy0opPKXCA6js
RIpYR3HID6qjzbz9MKTRU/LP5F9bz4pAUCNYCIWzkT8m9SQ8H42lGvTMsVOqsevRxCTSVg3QyWsS
oJr18W07BFveOeJp+LJfk+moM2gymBrT+KLwSfE39lVrAZFJI88ZX7ECJ42vMWBh7160jNL4zLbe
2Qm/ovL/3F+RrqipnHsA1a7qVdnpRZ8OAYm444FZlUlOfscZhSb/6puIZi5P4pfmfFdsGaL3QPbg
cjhniSU1Qwz5NPIFRbEfiwINnj86lywsn8r1+TMXXtC1cU1TwUC9pYxwnz6qwA1HQi98iIdJ1crM
MU+TCWCS6GS4TwuEnfx8heVoukRITKMFCVYmkRwJ17Jmi/vQDvg+shO7povmLjkL4Wd7ithAIAGr
98XT4iyzkvU+bEQTKcKTzZMaTWOj0SgStHX9MODHvtPdVro9RKmnveGRC7bmrdQfRredPkGlDdgO
WLzI4odoEwpZi5GDYiK8l68V31ili+Cjnm6LTaX0Z7HRJs61cEql0xKQ9ahKcUlU7DTmUVBqOwTF
YfHqIIffBWs4Hg8q9xQmKjMleF1Ap+bsAXW6jcP7gMS6oGvkCP0s/syrZwGgcdeJoU65cx6+sBmw
HUntk2YyExTz9tC/80BRt1n/oc4FhS8fs39WgzqOWYV8DOEwSN5ctt894Vu/1D2pFWiarVTkcgiT
ljdcTHbXQCoVvt2f3ER9RdKV5oO70eTxozzF2BtM1o5UVCk+obXzJKyOpi6sIDnRblaDKsluGwJm
3QHvrKp1BKFu8ZMmwijMS1Z70pcS+GyOeQOX3NQC7Fo5rhJR4FghaNp+Gu8nwkOpdHy+4rwLpiSJ
6u18PnqJx2O2mNEATHa/qr7N6YRESQ34SSj40vpO35BKdrtM6713LbBixBEQiY/qcfxH0XGZcovN
F8OJAHRybw5/8YquSZKw+MZg9pvH4YCBjGG/CqM70bvYLEHdWRzgm0Z7K6IhY2+ZCkJHPtAQjTuE
7w2m7Xs17u45eGKGm9o1ZTPN2oeJmT0AmyTNEHWczERb1rAf0gu8TVOKILjnCOne3W/hM9rpvyDP
hWesB1V9vcqMcB00jhiD2XtyI//+O+ew0mdBLzX5FUwbjBgDPYWx2lcL5A7PT/quFcHz2r38ggNW
JCN0FT1fH/Pzc+r8Sp3WTb28F1Rp19ymDz4r7YzPHEE61DipO3JLOGrROXP698/KQNajmvOCq+ax
Dmjre3di2KTgvLbC1A6QIY1lBO+3PLdOveSylF+GrevjqmKf2xmOiXZaxnhRiuqxGq2vxLKfEH7R
wK54SoDTNDxbE5X54+PDTwgdYHc6YpCiz2M8ikOF1arUn4zPtQXygAJJWUjWqDCB7gKbgZhL7572
m4kVeyM+vwKZFEaiLtQ3EZlCKiqGt1VqxX977f0eSnZyDYKrdhI8kwkJDSfyTnt+fyNDWmitASEP
Q2HIgU7RWCB03byOGh8tEo1NJWXw7WcvtKTekCy1d2wXdRAe6h32KViO0LiwWL1p7GG3kSrYD8i2
o/+08IJ7m9y2MWxO0JHHP+YroHDr8+pC+PIIAPNk9rfruczIpvHz0VhvS8NzbsqNahnuCMdV9se4
jpKByMwaDFGKfhHe/GaZSwJqoYSTC4OySHtUet8Fi0/TG/IcYOMUaJAA0B/npsv9Xwr7nCOQ2N35
FGvs73naJPNVqiTyZTr17WPaRHAe611ALRO9VorppAH8v3TBKXzbGliTVN7qwATDM+/e4soTcNIA
+/EwQ989LOYscOd3/bEZlFCjSxyMLJFPUiFnM7gYUxgqRQzNHZwH9gfIVacJ4WjMjDtFX5XNqoWH
R2DDaCkg0033UPsrb/hr/uhQ4ypoDCCQd1eE6DgMlG2YCMK2FSI7//0Zh5mPu2sFiDXWB3RQSA1O
kRZ6KEJSUrab7MWjEgpneIIv2RDoB2CfN4HvjMHjf0BH9d0F48aoCmSeQEezW7QUqgDBi3peqNb8
Hv44evrs3AwjyGSmBJcWJfH8DLDnQBxOFJZS+NgFdHV3yK5DQw56nAolcd0GrnTZHnIJ9zLyCjDT
vqZioZjXY6WDQrxFjSFq/r+gnDSY7/GF26OhhJicKimDyqI69WRvl5+P48SKRw1xw0HMkiou/uiu
7qyyJfzEP7+tVQ8tBS2VJUWq2amb8nuQnMWdt36Ev50F/NzFV0pQS6lMC/xQczh/ubnABQd7Avrp
gaSsxk87tUnbUAL1l9I5+fl7BcblYs4tzB7XAeYVidLDltJBZo8MTjdAD5x9IXrAwt8ENEd0OsK7
iuwxAN9ECOfjyyAzUPuxsktpL4nunT4PVFUypnJDVk6pIUlil3TgEDKcdHaet/P6ZpwamChzHoxn
q4IoKv9CZWy7VwpcPn/C3cZaR1GBitH1F3al68enCEfegnmma6vWFziyS0x+wgNp6GK4y20C02Mr
1Tq9uKN/bk3EHI9Cho15wBj3j5rzFMZpZY2J6lzXChkskbvGXGHGMjhhSNY+OTaao6CKbLwbTjuO
bRR6Rpt2u8nNvXGae4aLc1KA1DvGobKDuKjqdN8kYofZWDOi2PlbB/U4WrHd45eFfY3M5zzz5fWh
YyYTawoDQClVTeGZ7Cg/S5hoAVtH3rwsWxSAudB96I3SFUCWHGpvTWUbaw5MKDoMHpwigY/gZZlC
6b5IdrJG1VrTJyQOuGfhIl8nVYnHuYsIABu3ZPdxbvhUVS7si+reiWWUestriQR0MqilVHaGgXAB
fW7tRpoGi9c8uk/fQplZG7Nh5c4a/qL9HFOhHyVFLc2ZgQDol8cizek5rTHwKjZAFG+wz/WtqHl9
SGPrdpnnCpC1MqjAOEqxlbbVGIoVZ/Ub9AXdVh/FCRpPX9L2aCYZDKZd+f/o6hiKBoPt+Zvt7vps
sOm5L+eNfcYi1p0CJ88OSSFX6H5FxmNkda/p1OfMwA3U3X8+kd5m5gEogVhSXV/H9BASfAYRUDx2
pCstfOqxVBZ4B8wVhHDNheLGlVFcOQAOMEG036I13ylx8W+9brlKpDwwE6FUeQc4N2csKJqBjz5I
vdSC89MxNqiuTFm+e1CFFocTIe7gwxyG49O2it/YGz1WOb+S1BtLaP1GAmtLQZjBXCCirp9sXiq1
LNtdDJZsISZT8UxUUVGAjp/clRZN3eOSX0PPq1TD6jmSz9WNohUAWMZf7XJmChfzSb69HN5fEcnD
Qi5byS9T8ZxR14IfmcDvSikp7io8/31a6uxRluLwcXFFsrwTg4GyVussvBPVQcMHkNq85mwZqoyM
jGk1hpRmHw6xblxSofYui6s8BfbQleZVURI8vy5RkHWcK7kANnPF3btJxtBbvMOtRpM8w60/JYMM
B/0TaGIvYRC3CTncwaVG4dbf3f/VT0vsmJXkg3+VoIox/erfCSPR/XebPa5ng7ZVFsgg1vM4KflR
bKDlQ3H34olosqjOsLgxHh5W/p1wUw03RdHGupUVDfiy39fNVkd1gardXfIX1NaYm4sKLWrZzn/5
PJTBGeecrTbgNogH6bWOoJnqwNxAUuD7+uU24RCFFu0LN5qwTo+p3WP+CDx9twCECYsk1SbQVBpe
p8bs0d1jTSbRVbQ4RBhG83BxCmuqKLNMp9xwYAzTpnySrQWPIQMP1ECYnNEYdGP0XvZURLs4+ZEt
w3TzolFtVHUsEqkYO7Tgpl7kG5p2m5HWUAgDXH4npuzQBLZZo5eFZylLk6n0K83iM6Q9oejiEjrl
Y0akehaiayugq/zoixpM304tAiQq3MAmlWNWmy3TnydViPc648LJ4jqI2Jnwqu+OZetk3JEfGf19
8y1uSFAKTjMAu+AePWiiUw/yT7aAgVAdWqiKqX6JiNyc+/1y9oS+TEtIrSsn1aHGVq5PQ+xvG8bq
M2yMEr3Fbrh9SOY72zQCh2YsvSQIZuK0jkf26RwC+pPI9eRSxncx2ckFisHyZ0TB+8rU8xcj6edR
nYQUm2rFExwNkjGK7xaZJcdVEmXqqWJSyiJvxv615fMGBUQxOfdKlGBRPjQmE5MN1a+C2X6ls7/2
H0nFPFNfxepnSCzlj+Jhr5xCn2sRZM5kYPQ/xuJMtNK/epvCmx9kpt7cDGxooyLXaEUE/WUppnTq
X6z73eXbMlSLWjd5Z0AbKhRANTUr9cke+gtP0SJxk4QNStVc/ouGQu5dCAXMDunF7nD3PFEVqXl2
bd4FKtb8W7jXSCfWZzdyz38hfgAat8Sh7b+L2hVAgkIw3nYBYbfo6EdOOsVQfpZ5EYR7ar9cRRaF
u6yB0gEXO5QutSdJeqoZmW5J56hMfQrvJCKG+Jo6UPr+uBuHhjd1busdTI784+NPc0Zcbhu2+80L
RDtZ2zhOvbUjd9WFc2V30+mUIc3UyeEbH/DlN0KDX3RklIPNl2xxIH8H7dA8rzx0KeE7GfNIIoAR
JifZEPmbh/rk1IhcNFKmniDdpCbRSLNsXAGZvt27oP5/on59NoVAQn9V4R7yNCRt64n5B1cxTuRm
SLSJHHZSugYJLlg2JHWBNS75PkopV6d2pOc7xZd4Qm7IsMKLWnQVquRCfcFdAffTCIjJ9YfddRuP
TsWayApNGjgEVyDmply3WKQTqUxy3HDkqMZTJpxsr7Nbji8g+DatPwW3gEXoAfBwoK804Q9guUky
WSKRNDoTqurXMLgjAKy7zVnwRbiUW/GGrS6VaxMuzJlA9uIsm2YUCYQSj1VwDQzRFC6ZCBnc3Y8n
PEF9CqiS1S2YebgnIl4+NBSPsUUCeYMOtuGmzBj+DYmf9B8PES6r5jZzTPXZLUqjOQAVqC3kLC1L
la+1uqjPcsj1/Ti435z2kEH7jDpy2cpuvzkskho9ZldXzb2xpGMlmFD9ki1p9HNrSl7QNPjA+VKU
6hPUjOkNpYYAYv7D0pA0nwOhNFEA7ljK+OnRBr/eGTRLLlnZcP5gr3+82DgemX7wj8Fi4LvXRLN3
8NY4ZOiyaRJKWvYY0M/HhICX5e3/+r685K8H4h81SlFmr7J5WYHNFGb98bANoQJ1inYvw5CI1Iex
YMSb+ksnp3+8ynu9W7wKF5vl2PdEvwd8iXhGv9EfBknQsz0qEkoEjVfL98zurAl+AKwOQGKLrVlL
PsrTuXm0SOPucsjSiKaPYK5lIrXqvAgoUzqvhw7ztiXy3NsDTQBJlU0Zh/7mMCkKcHVJUjxdbSKo
iMr9TY0+pBPivtaUJ11lTQuAxM0XqxhkIl2BxHxs/N+1tqGf8oe0vxgmWnGhPunVkiYxrBQ8vFEg
9vu1ADAGFFrMp3LfJHdKC/7u0gk7KIPKXosU5s0zRhgc94E05rvNekAZxUt0nbpn8tr75mmaV1bB
ETdi8pfo0KS1da0UpWcnWuwsk2MWtw/pvuVP0rPaRnKLAbYqEO3feJlqpKlDOU94zhPb6LgduVis
8w9Sa3DNB3JjO58Zo+wwVLOScIyI6vlq90kLkA0m/pobgA1tfVd+qiYxsDzCZWcCp6dDXdFIi9+T
/x787wBeBTuzfmuyvtuLv7PvWJJ3tShc0u5CWERNAzO8L4/f9sDnzgzpSlk3JI+bF87Wzpv7cALn
uwv3yoFalh5kYjlehPhCdMKDE/lzspQJiuckLvnIoo4gVzVtlTA1c13t1IuMJbPFM+7yCCunWWVg
PWLVlqKq97n/Xy5aF76c6BM6LR/q6heR4nqPEpbc/0CZqBbz1StlO2bymp66Y4+MwlQ8e2OyvzXQ
VdjLk4WMH7sLa5GwSDVZCIsODSG5iZGF7dPeubiFdlqf7xzRHzc0D/q+evHDPD9AhU4MmOKj10i9
hutV16IgOaHe4dvBAm4rmW4pyby8IYJVwt24r20TggwkXVTl1Viker6G9gCAejRVUwUw9du+uFge
/sdqvMfpmwnEhVwNC1+q03SUlqi3U/2uOPJGwDJcNdeY07hIlLHHN5gDSZRL4ObIs7FdbzQMsvuV
aWdgs6vMxvcDYi5I6ZPZT9QXzz6I7y6g0bZX3uWsAJNJMajI1MnsWR+9YCnWUv5O259iWElrwKWo
IWDjgubMWn1Ld/7Cy/NZ33vdt2yUhk+DSJCAjkyFIn6OPIbxpUdwmsRE6gZfe3oYtf0vlA64e0fr
rsddDqv56MRN8bv9AfKfgXkRM30l//iWo1ElSf2bjEK+dD2Ds7964XsjE9E9blCwAW8bS0DXZFBX
iKBTEA63iO7DBQuyz4/r5VGPkr75iKCbF6sNgK2MK15PhKP62JIyI9TrKcVJwYfn8VUSi54cYmkz
miosixA9PVT1s5HtazJm0AYs4EyrxqE9Op/zVu5s0roXEqGdmhzwdCMFZF83coqWsEwg91o8IXT5
MrEK2jO3GSHkxUe/vx4DfH3XvqECcPYoZqivsoUDgLHXv5nzFE3o1rCSCXeYmwDbVX5Osnba9Q/9
lr8sJneVpZ+IbGJ5ktwKCyxyFTsDPc9C/Fbk/HwwSC5UFoIOVkBzS7+KeQgdHz7Pk3ppIMj+BgoL
bplWj0PK+L+qx72lloElSaVl0k/mR1NtWQnCZmLOIu14BZTQi3olqhVV+t2M1fQDwi7vJKnCFfsN
MiJOAHS3TlREo7PQ0XZLGohy83+EeRWF/Vojtb8S64l39cy184W4FGK/inEi26epwj1lbbaEFDN8
hBeeviXX3ejX+/iyL7tMrNCmiPhrwHiCBIi5rv6sqVahxovk1QcIj204Nb37tFC2gs3Sy7EW2zq7
KecZLaEw9aGLKYYyW7j0xXe0LsimlhYO709FuSEBaV6RjnLIeJlaJDu3E/fubgZmMVHdXBp+9sv2
F+CvfVPromzAMfBsqj7S6FBp2d9W/T1MaYT7t9LD+IcPXp3SD3TwDfi558U4e7AgDcXW2A5v6nxv
HxQLMWYMIY7DTq2zJn/6VdA6B31F+kvNbxAZ1jfGEMH95xeAhh1QjJ45it9PogzBC1xTBlvIAj50
SYcoVb2447tyLgyhWFd9zMnppztN7jNvNkvP762vSwO3wgMHSa/dbYUpRYaSmFweIYH5vMN9hy8+
UH9eAs3CZQr1M7CLqNE4eQuaWX8PCZ7SJm0EMVp650u7t7s/na6S1K/Z3rL1FOisvcXbhPJNsChz
dTr47a0mqMfOOGm3hFPGzy5ZFMNfd0dBlt181bff8P32tMAD6oX617xCIgJ0X0p0TicX0O2p1W0P
wbjR5Loh+LhNUd29SpUyj/YNixneuR2vlsMRNv+WcVkmiP+QRSR8cKPGWit+zLA2ON9OO8H0VdWH
j2Ihvbw0NxxIjsi1R4Q4AV1mU7ghv4llM8BmeF16H6Ber8AZpwY9h9zbxJAuGSM4xGXgyfqMwKRF
HhNtqJwZBnoc+g6ZLtXMmye75w+tiXgFdySdqrDc3UfDezoUErPbHK61GCYYffCfq4hqNObACM4q
KS5vN7qdLa/wDmwFxtZMCUcSoKIyv6VbNXg/EwJjUQr0I1jBO5KgsxQoiDtPSZA3TTiuH1z4jlNe
ubCuC5ED47xeEeznxH36uLy+p5uNVoSkMOXoN8GDp1iOlTZHFZuWlJQrtXXX+BITac2MrZrq57Eu
0I20j+3Qu09iWqzU6SD4byaD5iQ/w/YbgE2F3zNSHl3s6OYI6hU7fcrNb4XS6GAhK+HFi7BddhTc
Ohfeks59/ICoAWqmpE9c7GO1Sd2f9i/4A2NDHjz64rIcfSv1EouVxyp7HsKJ/nBZAk77Bkokdu3r
zlK47YZl10kBiYTQHck1mA+MauQAh9ZeudIp4CZNKt+BI63vfH+oFTYpSvysFNBF2ZMP4aytufzi
A/rAaJK6JfwugTOqU82va3o6eU5brIu2TEWMdgWD8hTrDBw599uxj0kyKtXswJhGAlCdqfmWATKf
uBzvWMr9AflAA/qK1jhRBLuA36TpVIKYqSWS3gnst9koXDopQN8VFIuNiFhBzNGX2/dXGf0Ommzs
kF/+qIa4POU+Gr03UAbPB1cRFeCIR7XggFq5hwKnZ3dLYicDmIiFDUU8Ea2gbgPlaipvLbzvxycv
9TPPxsrm4qCmvgbvdCOYjHE19j23zhiH371smeoTkAQ22IBIuwg5tHY1qjiNs5+cRCbYC5DsJI+X
T/MnYecKcEP93DDavGCPCshGQOU4lVEexcrpRre2lr6nEtJFfUBDl1jxgMZuEbr2JUaQs3QoGfTZ
cxbgJXAj/LZN3sJoTRj+TKG2j312BjxbzGanun3EctvH9Db9d/9JpR6RMOCCLkt1mA1B3M8Cq+Mn
Rw09FiO/4HZ/Yq3Zs2/tkCr/FmR1VeQ10mybLcDy7rubZGLx3m58jciEZdM08Phb/BMnCwN953VS
ZDHDYjQtzdw1TjALY8OMYYjt1KMFbVQB9+sNSzaVBJa0MDBwlv/BbV3IB5bmO8xBkzzBe9tJ16gT
CY5Qz/tjmLf5ZrtOF4h0Cy8uCw3E+p/T4Fs5CF6mYuTbn7ZIPv55famnsX6v79Mbx9QoPLKBqB8S
TJs/2zwKVKvMPGHKBf4Ds329tkflrhmQN3Ah0KNb2BTJxStk8Q1JsHdTYCgq5wIzaQLspMntr7Ls
H1d/cXtauM+ewXCzrKYX/+3tEXrfb6t2J9PRIvZD/c++mw8RGAUUKyIVlj+BY41npkMfTPdSk/gx
0j0qgMEvmT/OnD9ilI7cJt4QNvbSv/NRG3N74eh1vpnjN+hkekqur2va2hXMHdv2qdbtKQWIeuS4
ieCvaQcwxhpZ3uliTqUgMf+wN7NdCoIoWPG+cmBdbDc7hyhvjVu9gmCJKcdIW1thiZfHaQQwBEDj
22fEXkRcevO8qL67o3vWkY1Je305LLn/0C6UIewLtbJO1BvOaH6DZEao4pHvHgwzi/OcITSYW6iI
KpvXmRqq12Lr+i605ymlL9mowiUur7KNbs3GaQ1VmGCNfQtLs1V5iCPD9dtDkwi5Q2HhY0gwPDBQ
GTmluHdtr4/QUZl7gy51XqJAvEZy0pVe0KIJlJLKLvXQDFNk0EPpl8n6aWpAiZwxsn+jSZ0UFWd8
VYn6r+MqqS5BbPate/dwfB+Dzy67XrvTOIV9ZbkEnqfQhviu8zYBMFWzf85UioE3AdfJmCNyoGC3
gW3AyXdIOJkDuuhdPd8uA7ilY3JZGg3COlQVLhsDAiLqW+xfMyrlYijZ344ZlqIJ9BkYbMZthlFC
ew0oPOATOsSck8yHfS7r/DfCCG/wOm8hMR/u5fDNS503nphPI/SjiIcm0P/dIBVKgc5mFfbV6G7q
w2izNtfzDOHhfdwl1uprRJi4GGWkrqKDrlO3ytyrspeWod3Gf5WO8wcXhq9pE7G1ICKfxUJBVhTZ
Rzgn3l8Ya7jGjdQtTacUz9kYGCIPcpl6eh6nFOBBJ+T7zT4eZ6KwFMkK1zqwVnxKmrONLUxtJ5H+
972l7EafORVGJnEJnqHDbe97xK8FxqMB85S1CyVVj6QYAqbZ3zfh+epd5XlMtlWehLOYLOoAQgwm
P1uWb4gHdHu5ymfFjhauiJg7wxYjXMYOV7QEH2GhZ9mjYhLibf2DvbbFL23XVWrJPfDZxVaeSRtG
FqRxAUO5Cr3tIVCF+D3scaIzNPDcrHS8kLqG8lK1iDXwFSYexu9mIuRD0ghleGID8o6pdyiDG3Cx
PGtOgISWcEVpvNT/aZKUQa5I9oDD1fZdtVdiyyaCFgv8DVVgxLkggjNEncL8+nLaIv0qhl2h781G
aWMcpOvi3Qwv7jy5ZGp4RnPH5uOoDF6XwVnk6Gsnwp6c6mv7iEN/qIF9EImOsKpDDjhHLftgJO61
5o//YVTDnBAyfHXLtNN7WOs2JW3x79bekleApi7xCyTJnCR7QhOhuAeBwLr2VBWEYliFxAwmnIdb
YsboWBjHNDn2Pt3jTda6AQdL2n987laZW1CakzSDzkMzMSOgF1w8K7FNzYcqsVrG8WVyEKCIrrET
LzNRw1B9jB/5xX0iNcRNjVtkj0QA5Y3oJLdFhPXES78/c6Q1aqkIlsCEIFChFXjZsWCVpagMR/uM
iwxfA4weQzwNabueK/7V7IioGXjOktSJLkFru6zag0Gz2Yt5P7p/rgqxQpDmRjNDRzjxQeYPrqWO
d7oiOQMdt0YMa5HCZ/khBGnEjU1ozrplsNwhgdM1ZkE98r0mVz4Z+5519oWySNCoKVoeUFELX/Z/
JGHaiJVBwfQtgXMNS+XWLyKKDJly0/VjETuLKhsqgep/LE8+atiQ5NbMrCLlINuoAuE2unOlVbmT
ONS685gdh7uWwSisFbi9t68qkn7v8u4q34Wo4xL6FfUi5DUs0dtNms+I6AlcPUEQsRCidpRNRCMJ
Fpxg5fqXUYygxQ8mjNwRNR1VVOTM99K42eYMQYy3TuKlXfH4L1+usqh3i0r/yiXoABi2npL9WIz0
1pp4z3Ov1bZHqkpjUGBLvCXPV6UjJ2nSouSodl7VQohRFxoj3YUDyznLLV0RuybKjB/0Sd+hxDKn
GevqE8UiiA8aun/uQsuQmVUmqMUqf9qioouEfgX8Xn8l848U/cujjRg+5PI6Fc0povTFnVzIYjnf
8sR15Zg5KqiSKO+9fHd4NgO+T0imEt16mtVPrWlN09fp/LwTNmRetcnZjdAn7Ivx+30Vz1koOdbq
hCd/hFGomj0MEvjJhCU5J6pTeNtB14oxWZcBFvf1p1rZlZZvZGwGzIQ5wvzlH34z9Ib9SvWSVUWo
iCfk9ORhJR6K0CkL2KgWBz0acsM2Qbb54e7dJIp0v/ejM3wCmD/Ound1CkeCKxO8oLDDuRpo0zGY
QzggURBP1j7of/ipw7WB3ynvyfw/k/GBBomEWlNQzyIr9evj8+eVHCI+KaAd+gTBmUK+m8q2BVeH
w/95WdaRlGJYjJH4WY6JOG2atCbzJwf1gyJfQ19FB/6XVaGpJj8g8ACatnU7TXwYOh5ipuxUKACb
rf8rr9342NzQQXS2RiAVUTfjcVL97vogI72lr7Si3nh15dnLd8YWQJdst/xWeMcUaK7XPe3Tlmu4
3nEKuetFAo61Bw2E+jw7AL1QJvyVNBNXcLYb8nYHXEHezyUxpYo8FUCYCSUC2nXMfGmGRepq70MX
yTjztaeCAI9l4sX63u0vlWbev1Akf+x7+w7n5OiZ0QBlyXqnQZxilMtmNfJwS8DOCCvgKhwX+5yu
Ki8MGxoOn5Z+z6hx01Kj+6z7Mg765cPBNh5z2wGqUBMYMx1fkjYgoQgEwmvo7lNJjBfvM/mKl77/
/bJWOXVWwo+Wy5u3vQtexgofgpuP/53SEuY/R8Qdrmmtq7EzAXkP001LzaTm7GUJI4JKnK85x2QY
xzZwHlQ+l/tz3H7zMCeung6EqD6+hVl0+bbL+12LNOpqHf6OxzB7FzfbXvn/hgzUdizZRWykUTRZ
Wi0W+uuRqrfRnYYNVNnA1JLfRd8iRAAJt57U9Ij6DfXVdFv0rRp4PL74Q7n47BJ/JaDqbuKo7QB3
R6TldUSr5QXKPPi1HeVCCJudDSjU5sY/eInX5479EZrCYsAFJygyk4o6hpCTK/kX7Mgj63+mWvld
gIEWlMeuwcHhDpX4jh9JqE3G775arF357eVCsOlTykcfnpD8AQ0l1pcrFBtkbOhpRx3xbsfCpuzz
SKdGE5obY1YCR8/JNoCu9OwCRw0ZqelA0eczhSFj3aDy8BEVsCtLX/2n56jFypOqlN6pKmWHRAxW
41DW77Yb8BZecUeyr6K4uEsCTlpGkzX2VCyubHIzpjkcIql5saCDdDIdh/YA7woD1qWdjMJP3P/a
DLr1RYgIi9p6eInD7NiWQallgHKzQrZqWjzVwYsg4Mj2pavHw/WYpymGpUoLd50DlZJO9ITbJ0wA
kBbJI4bJB9mxWcocaQUQUfFOlj4C7BSil+apQ6h+1JWIZFHVHlzL46qpYR7DSfjHKO2xKa5H0E1y
6jiYnDUSZmZV6g4jNT1y8mHuuEIrCuhhrO2iiTmuR8dr32FgpDD4eX6h5oWWK0oKE7KqCYQp/amP
5NfABqfXO3YaTDX9ij2RsljYqLgTuWeueDeZf/yutWdDo0JH0hdhdSxgMNHaAVoCzD3Bi+UwkyPW
GJ3+aMo/wchl+Aor5KeVxJy5Z92dsYpLX8xiLDBnGqWQFtrji+qWUNvGJp3nvdp+zD7wqsqBjb3+
/JFAAJCLe/X5ei7WkxjVTPS5ng3V5AMDQi3Ag4pa7htkHH+xyCBlnJ23ppOefB0D3Twcd3qMbTXm
B/CpoevaRfmvv6m84AVUocXIBKhHpVvfJ3d4kErJWUGigGxstwz1WhPkMnzHmHKP/0f58vESxbve
XLs7QSkRxjjQYVW5kpG1oOGLv1WtuSyapU0LvoivmUe2Kk2mBfUX2msXl8E8I7ncyOyabGSLtReL
KXrk6as/axhkV9P328iU2YQZL3PnM4oP21sAFlF4GmCXkZ+LLnx3Ui388cxkBrEYHe7pgCeKe6mw
lk+BsRYiEK/bT6flN+nLWqgr5vf69kyEVrQ5Z0ZRPwow6PTOzWZMQ6+yI6Lwe0E8MPxkiUQneNQX
/ecyQu20/v2jLjdNmQhSUOnDgxMbnxakudbEiDMXnKc/6oZZOa0iagfSfinTDkS8pBJWbliOd5UP
9GheZekvWfH6Qzgxk7vqwXxjaM/w5ReuHFFWWfuFv4dMhaNSBoJ4rUX0g77OuRl9MeOK1NKuaE2r
KQ62GL3gLjboo4+3RQXDxBqYYS33pyhhpvZraqOH9DinDEgJNJyFBNFzSwDfgGrex4tUcLKrIPIX
ZnGn8GdfxepVdVVdW77qw33F268KDJtCw0Xa1yJgqi8epo8CrOSIcFwDFGGh4AprKKbTuscMu0AJ
kXRE1rnfls7jZv6RYPkFpPHEPESg1VonJuO0yE/BWCj7CumEOHr2wpnYBFbfNz/wo6i9qBMUJl8m
ZluvBToMmIUGNCkSgfI2eu1CM4Z7lxieyid3CIbYMy8mUhxkkILK3chDSA4ONNwCNXug01tvO0TU
jRNcoSTHgsyZZ7yBcLupLzcWRfOX57B+0nnlRjTlIALz6QpvGA4AGr/nE+3BDZmQRprVVg8xifaf
mjXet0Lzp/hmrmoQWgSdTQdZJDijT04SbAImIKu0by9svbtpP0dipqbA4yRUaCo0uyiiXMA543YK
1mXf3A3A0s3oOEZO+RDba+qmJ6NSdnM3wRnZEWrGiSN85jaChHyed2vVue6MUM+EOesZxxQtSkQQ
8gr1dXs8ENDnt7MRs6uJPBxCgnAWPlnYEpsV8ogKElQ8RpwGZpYQKAcm/HcD9Wzhm4Q4tFYEgu2b
bARxMtTT5KwwfbmpkF2k/BFv51/QoZcnEwE5DDNsNsIHiR0KMUQVI7c6i3+IPTkJebjRwsegDW6X
+FHRDsz96MwiRGgBaYFCYMwBpqFPcWv/RDhbr9RqiChxKjZXzpqTpkoLk3N32z+/hwndFYvPdtzK
6rvKKQhIIS/CPAvVec9LnAZ420+hm+nDR9ehvUUJKIZCUK3Vz3Z6wDPcTAGcQsdBTJ6PzUv46sFw
GZ1XUEvRraWp/RIT8JuI2oyCUVKr0dSYpQjxDlQCNux6SG4Si7pGMkjVsNJ8yo/iNULC7B4GeKa8
dxEmkHWJQi6Q/XaKaFgSUH6wGSeboJYqYjREzZOuZQrmK0ykuPgEEdWnqtbcfpJNLasF0oFaP9Qo
9n7LaNzOWcQuKYpxY1OckoVKoQzIW1RxTWwyDmO9+MVwSIJsaLcA6LKYRp4eFPjjpAhTKEUiaz14
BO9vJtQhaVmZcUx8Hw3oDseG79Eyq40jHNYV/hwVymaw/qBBQcyKq7gf9f7OodUK0dxZ+9fzBlWW
QTD95R+h3nymIxx6t5iZminO5geLQpVCHEf4/01296SvE3WrCwJlGF+Ys+hMyEjNEKRoCD8cK+9f
GiqvbMmkmjf5UtEPTbbUTRzNJ/1b7FAFERbMyuyPmuUIU1nh1FtVIijxpqRzOYgU9c3/gM8soDBu
tes445POXoYata/KT+K0YI+ugwb1b1xgvAAYbcEZe4N0w8vVI4JSwwMOpeeaikGu/e2Lky4JaS6a
jhoNHxBoNXctnzLGHECN4vWnpTMSL/gpoaUVV7W14DNr38Adx+Hy7oegID13YBb+Mddm2iWI1kgP
oCfj880H7yehE80+8Hhaf6OjZgIo+5FVbp3966Ki8jodFRjkVHu4m6zuXDxc7zufRC7UwTA1o/Vq
nTjbI6LDkZBvT2Q8pWsm7ZMDUsYUZsXZG7dARGciFkWU64SUSFkbAVuXi4Y/s68qTIm9nnk+BrHW
uq8hmhKppuncnjsiT2FcF7BIMsxe0Ablsj31D4qA03CVYBq9X8gc9fu4ia2S1tIZ5gb/ndTyl8Ty
Q5ULSYm9Oow4hQa6qjuKdzms8q2p7/VGQEi3ErX0sQq7TW7fHcklEhVy/+TwCBB0OyPR9nSxT9H1
Js3dVcPG7CBJDb1o0TXdlKm9lWMyc8A17EKofBuu0maCmNUP489VnMlynsX2bFLtxAREPGcKaC/E
6r50vBuKQiFisBScFhhRToiJATZ3LiC1xq7dl14e9G3wbd27kzlpqYxUluN2mBphpok8iclnEi2Z
nJjCrYtdDx3tLAcPTFhE4fbtlF35N8Q3te5OPmlgU6JqFH7Ir+FVTYyzerlZ1+04xBuIXkKYFoQh
f92tSiMHoVhS9vIm9CM08VRb/rhl603SFHgwEbYdG81ZWfOOpP6hKWJ9HfQD6uSUwh8xNcHRdZiE
4kinHKOVm/VUYfShkl/oJK11YSCXMU1Slpww7Jq+uHmpVNC+94kv56tIgLlpZtcIAcmcHYMYiF8R
4jzetcWxv+oUsDMUyI7G26StAHGPs9XsNTNllCEV5AAllTwdfzHAZsFpVn6j/GFicJprTmGBSHhh
9jGZ5b1MOJocum2VDI7ngSJfse3AWQu0IU5v0DkmgAgp8akKZbrInXRGiJ5PDjXZhcpi/WvXeFwR
ZNrAtOv+aG1B/X3FioS7kXix9zatFZDBTh14uXLbUNnWqbusrfyQuBT5ZAjUz+iXrhRt7NdTx85b
hwpPApzRQsqSch7aRWmDI6M6ZYKoDONnSWOrFkGm2HKPvPq/w+z5WFX/HTOsaGqNy540qkG47B+b
aVm2n4tmXtoVrDcMXhZBI2568pD3u5Ik3q3wNzo7zGp9qLxocD0ShyKJkX7PlyRUSBDonDAmUKRW
++dFdr5UOKX89JnkonQ9H8N1RaJdgdv39s0uZDc44C2oGfMSbl2jCc0jM+ttXikF8dUfNrCuy+uy
4Vyod9DJR0HZBpeN4h/MyTSYXcNrRjdUTUjtXZG2Etir6eydvbhRP+CzJjgkL3QbxLiv4+Ldnzb9
f6YZw3J3rQ2AgDWkSc76x2tUOwvUjm82XBrbAFxW7/hwKCtcw+IclMk51vZO2WuiS8i7eBYpPwg9
zgojfSTqwP3XGg4Ej1FbXJqhaQKd0zefE5i/ojnPLgGPs7/6SG53R+zdNyF20ru8NHRG9kplaw3r
M5gNM/IatP9q6wKJ/gzIfTNuPdO8pKlck3JwfK/2OTCQ3L2tU0pwllc5olUM3+alhmvxSdcZSJmT
C1sWEr/sENbiO9kSKaGnl0M5D0Aob4Ba7+iuEVhwYtOLi08XnAqRf+I3/n5ZEqmoiF4FwkEs51mU
7XTF5r079jRkaKh+ERP9RHX9RPfpfaZ9MdFxzXv+hJm5+xGPrblH2c/FnLKRq30G2RlBETfhznpZ
WVqOgmtUbdzBqpaM/Lh6ync+Joh1b2lK1bqVXFb7oPJbHuwxnHmMPBoU1DcC48jQZWAmIiXRt79A
pzYmDmYxPZn/KS1tLnTAgWybb8hUfLuyApML6AaevHjeZOddXtLSYXBebr2UJIl2qWtU6ZXlYsDU
/Bshd+EnNfMYbCEpYNmkdOLnUra5YlRIozARDaF4934JKYt77tqX+2982JBZxngPZN/AJXgQ3zpT
X/cyjNEjs4T/rT4I98exuixGiGx1UYH5FOLQ+qHkg4vutvddtl4VjjbYGYXS2cfSt8q9MHGbK01D
vO+0qdAFTd6Gv02X7SUjsvFG0qICxDKU41Q6ql4Z4ZnrDj4r97Esgqakio+jGTLbAPaJCOV+fV9D
RjUXpHU88vKKTxNBnHoKk/hRsxBZfm2VhmugKvIQ4GNA6+UHKCFWimHrnQFthdI4H8kxq3NS5Y9L
FkLNhiclg2pCrTH8VESvTUI8kDCxDOMrCpGVdzl0G2cIC1ibTNDP2nt8ebmn6o22DcuEBOXm6wMX
tDdB4e3GLPfI5wTGSH3chZay5PDaVtbN7pHiQ+CBJxtcP7zFppLovGAsEw9+5O9HdkS7YBzWflZs
ZnNPHLK+GRhXEDx+uUtTSlTg3SskEFCvabDcBj4G48fKk/B1q+xkLVmW2UOs6gBhoMGCH4Qnac0Q
jXwlYBCHUuvWvO4QV9yLQP3uH7xLPKZOlZevcuTPgRjmmL5sacp6kac2VYo76Xgsnsi5gWvLZVCt
RchjHH1+1JqK+i/RLH/Ri2ZDRW4UB5Om/7jRR406MqAQmbPoccuf8Otb65np+IRetadU69AyEvhM
2DvFn85MUHJt46y9ebuGg38gFWOziSytySJkRl6FI/qkwn2r1JflJsiPXb6PYjISPPfTuRwbe4pY
uUKmn4BZiCE52CD65rNuKBoXCweP0QsRo1bb+JaaWxKdwPqma3/gAc3toAIk1g+qR/PXnmzHGrJE
T6oRLs19/8hdiyj0eKmvQTnCuVMgBw4UmCsT7SjU0nGrww8dD+j8MseCFjHzRtXyae6X0DgBBMTc
jmKjvJsyDI+Ncmbvjy3EGYty6cXbZ5NbkGoAHNBDzYKAeAq2y+xYFcp5AErNe3/TH37wnKyQJBUh
KUvv0SP7mOZ57cHFI9l184klc8a4wsYbBElE1Ex4MnINbY3ALwHu8jSIA4QxjtkNt1Wu0gvwFD+/
8K0qiCyzrVTlvUzyP/JnvydmpROcwFP4AK9+ge/k5y70hxmdxDseSbKUaPuHh3haH1Bt62ppLpoz
RFSmynGB/+/PlptzKUmKvY851T4N38gPqmaWDCE3BGnXj/QAgT3jHjkuiM41hkKX+yT3/6EzDBDO
X/xHxjeJuqwkBeBfYJXpDdP+llnSApTcuq0Klq6l7uBPUpcxZljt56QDJkEQJ40zscTsIUaIYCKR
mB4rT4gQCSgTmc+PTe2tWxohyyG6dtOkS/JKE1pF7tTQYFfgdCh6ZpVD+YRMkImRvC79/YPt3abl
kVH1MLGil+x2ZM8+ujuBhKrsOZHcgdiNJ4YlJMUYCt+djwOZ05yJ+Ay06eS021Yq3QMZsrGaJ1bO
cr36s5plhN/yb+t0PA96q2IyTwzV9dn578PD5udZgd8CW8n4ScJKvsregvy3cIeE0FytDzRkgpkv
ZLC6MNt7z9Qv0BQAdMHk3GQCz+KbcnwP1nwvVIRDo2nxfonDJd1qcK9qWnaRmCeFp9eN6CEop7T/
o/e7X4cjGd20ePuLCscWY9Og0p8DokgeEGYwTKj/XsveBBzuReYuPY/7sw3cjULGZTDeTW08Tbve
Gv6+nDDKaphu8HAMXeAKHHgqSOJSPiNZk3OHFLdlX3xhR4s4z+SHvgwpxUcsy91CfqNvSsi1V2Wj
g3m7PJtGkVDmhvWCelfjecvtWEe+rhNWSfjFqh60Whf8IYLQai63sryvnTR7NAcv6sgT4a2Y4Fif
Pc+sM/eTu8rWq1woS46hZVqLzeVgeZCTjsckfRbdlZxLPr3I19VFr2ljX7FPfQ9D16Ch892eMErB
c6cKCVuO/BJJ88ZXHvKuY5y4wh2NRhO/naOvQUNJpIK+QcPLKtbsp7dZbI3SwHmZmNtCz8tQngJO
7ziGHUoXxroL14+b+Q02n9FsTarta1cvZmVY+R0X/C2ISCJuGxM+m5tJUX+Gf4T5MXEnVMg9pxdN
9LDDoKV0UzslIQAbI3kXOh3MAgyke7dwFKdPgv7mrlz+jk/gN7zEq9EDiAQjvuS8kb08pBb5vExo
jYwJQX8p3KaUwbUJEW3qenVpn8OJ24GEa+O4C6nQ3YFkoIudnRch71KEnAKDdIfNKV1ieUtyFgox
2XMW2CshoDPzorLIfrWoIwTpX9n1vhxjnzBisyQuloSaffSQGBxowxcTdEVwWnpT5KgCqTLld2qR
47rKFxj6or/anNUxsTGYPqwawESlIUYwVGaD7gtqriAozW9EHpocgs2fplw0dgqtJ2kPmCf6JEL0
sM6Mi943vlJe5K79iBcrfwlsB1HL+DmVlLMkaw6zr8X36sY3PROZECx5KXwY9VBmm+GPxAn+NUUw
G6L0UQODELqfHdQEs4w7LtyRFfUbNhSJKFZxBfKCA49tnQ/rJQOsHl/CrIrtC8cSKcor4ocPExKO
WdptndfCw6oAokNWjrpEfD/iQz5dqn4i3y1AfsgG2pjhB6P1enRlIIg0QkhgVqfeXaBo9uUQbZCJ
qTCGaAemyRmnsv5yF74gClgCtVfsnvcpRx9g3ApQw2tVHggEPsnH1kvAsvzp0A4R9cygc2XPAU2T
iqLp1d14o3h4mP8y/Pyuz4iEl+rSa3P1SLxI2R2RMljCfxmasegrRiiSGttDaoDMIXn9N4zzlh0B
zLhpYPaE5W0IwV5aF+cksauPlH9PDsjWbT/Jr+gbN8vOZWFHdZ2CM7mxNubIy8tKUSccmETnGEHz
rneZSEn+kmoumyLifSqzhmaDbT8cw2693vr+UK7BIOEjEBAB6kM/hTolEFAOimdRbc6XRsYgtcAp
wT7t4p5l6T2DnlvxBMEigxD7sDqpy1rMG2yZ3AXIzJb8wCfCVBEJLOMyWk4lUHsfX4W2cwJD/c8+
qDsiVsMrJLy7K9HyL/CZuOUFVY2oWumh418VL7FlKV/+AeZT0/GGbV/SxMztewfx+YkKui6ZcuoO
ZnSmG55nCp9oqqqS0nM5ujRy6c7kTH/lbwFOVXJgC+8f2VKQqiJjha85djIKK+1HEte7JSlGazb5
ihthZjd89zCOiAkrlu6MLtsLbW0M/E+KnWMbnwpFMe1fRhBM4EMGhr+GhRuh22DM46sxBPk19JgJ
PkiH0D4XpCOG8GjWJ+R8vdzDM/1Xeve0OztpDou8gorW7+J5hl8i6RKfrEtOAgRXjH6/2tAg7+Yy
3fkV5itilbzXUlV3qj5RGWV2ai32aFSnyDzUczlWRjRSi56czxcHNihTS6wnRjcSU+XVpcftFRP5
0uR3UV49BOBw7MtOMn50amTsk+epA/faxO+Rk7TlAnO+XazTNThp65iTZvlGn9fKgN4zbt5mMqSY
GAxCRHufotdBwVOZbkzToOGsJDZXV4n6KMRe08cVmjaI12F8Hhx3KX6Zix6q+wx12dU4IL3wM3nX
3P9TPOPLp1+PV0Zlouim+ZWSP8MR6xbj/3zmL8p4mjvWNMj+fQyhKRsbwRI/b7h9/qttm/nEuNiw
qGm+gqWWTioXkgN17H5LO5FdAyk3gyhlySDOgMYsvvWOzXGtKvIEKiex2gU48i14hxEKfjTuxlIh
kA2PbjYXBORpRG6fbAYcu/6jmG8egLxfLknC1HChcU+PHN/WBx+2GflUWDcEAt/SwO3duBcLRAAc
JsFIh8uDqIB8r2qM9PUAWkyjDK3FlVjZpM5uY0W3kSmmVYVrKxf6MkVcRI62VxB9EW9oTTSQoWwB
CPxnZ0rCufDj6Cb/dNwDSa1/RnpgzqvjYPz22lq4sKOxkc662BqatB6jVQsnMwqRTsi0Zq9XGNyQ
4Dj8dQRhwbC64ONOPL1TqwN2Ob4iKqEs7vRzB2M0OVvIaRt/01PT8cHcuE4It81gfiM2EUaIgrZ9
NEh9c+5eCyeXxKFDUC9q2POT6I8ocB+7A8rAFhqdewdlA569dQYwwbx5QdUCuzuCxwZYWxNiGhJq
kdJb1R4vFoA7+MhoesvtNuc/3+Oyb0Tug7mz9uRRgJjS8TngNaG4ZQ2nZY0eBAF6kZQ37vYh/Y5c
3t3lAlunD8ywlRm7xLHl3/fvsRqFQJt08NnPx3p2108weRQUOQkwwBTxLTPq+bzmkjwBigUPgTJY
Q3MkdlhpgDEN5HwpBptMvVWW3J2tQhPw4HbHHz1VF+QtNPDnos2cRRZK0Nu7mqrdwTu74IE4iLpT
QbWPcdBP1SE5IyCOIjU/Qve0Doe+yVnV7Q5wNbABrGMLuzGxAiqsz6mEivaRfL3TbGMhl71lMV0K
5fo3gQweiPWX8BEtISovc40cyy8/XWUs86zjrXVowJGwvdwtkDVKkVUv/lwuWFtXnBGeZ6tM0whP
0A/oGasn9uxSxELQZmOrqU5xHkc3+fx8gWyMrFpdozNJ3VP53Idgkh4ANk/NrOIG2yDRpxb1EK48
DFk76NPdYQPcoodQQG6n3MBGn9ZPJDiyRRrfFBWvpb7J8I7wmtRgJ2nzn8bof44UVmkhgRkXMlhE
sO0xRTavu1g+DV5fOjVmKVQfnPEsr7aqA85QB46mCGNSLWO2U3tyU6BGN48ZwToBQxQZQcbwdiRI
ZVZlUI4rlDFRzdTbbCSlF71KWFuR/23+BOPjYUbcLrc7GlOiPq1MvtQIaojzPsiw3aOfN6VOKHeC
6vM8sbbf2s/RDOlH7ooebHIJRPb6ml8TwBbif0AV7dKBUj3xxPbfjWV9UAc6Ajko3OPIbGwdFGkO
hWuxHJCNORRYjtGtIEXJsxnMwXqhJPnFsV+qIrapjXy09YuZoYTfXuWi7DxAOtoWuTGwjB0rtDwI
NNkluX1ZKDZkh9r3vJA6URemaO7ibFXolt7cO81BOaspn2bgj3VLXlRGMNbXmEboWe+sowFEYYCx
LjNGy9/pow0Pf4gp5A09k+lKnQSuA9f1zqdeeQ5X4YvUA6m4Tg5QFMT+YdssByMzfTuhII+Isy2c
2si5iFEjIe50JlfdJRlknClAg8cMsN1QW8N50quWKwLcn2GEF26ozimAMQ+NqcTyLxXTwJV0gfoP
NvjJK1zcc461f57qHEiEy31tqwxvt4gi3rvekJNX5HilNxCrgnq0vI11s2TuLW/ZzDUlNArBOzVe
AvMbEmb6/RAzVadd8uXf/00g1j3wqv+Eu7KqtEFrTm+4OyrRkKahktMm3xDfUuIQGnyDrgPUx5Km
M3u3onYSwTSFkUjmCyYmySkTJUucVwe0fP+nnHYr3NigUsPhxauJSwsrQrCVYZs2MP5fqplze1Y0
8FBHZToXCHXAzqobKjChkBV3h2jw0t5zgnlblKZP2/BTNRVZetDtij0anSGM6GukHV02X+qTgFpz
Vsct9UgMCy9olvhQ6hzrQIZs2PvnChJcajJbT0DAq6jU9ze8ugQcfaJ1oJ1IsjlpWrhFHO8PIGmn
hqtEU+Ra4Y+fMFDBZ8Ew8pLpwnDPpMyOupRer0tpUriA+wc5d7AOT5/mkEEtILvIqeyTnyGac6JB
9SvYOv/+7fZW++pLQevsXYjJwyJSFAQUSY/9tSbhouccnGm5xgVXiOQ1tfMs6z7PWjAfo0vKTAZY
5eLNakCeQDlKhV/SL8FqDQ5BxR5fRba7xc/dEb4c0at60FOSKnB2NW1HDZqyiPH5IftMxZ4lIAVD
YWJ+hdNAj5k611jShhiV8rVbqF7vsQgiixVXZKRJAbniPS0+g62tozG2/x4JgkTyiAmJRFu0CXsM
imCxcz5ovWDtZojT9a+qQ+iNkHNIViqIOGDYAxljMmuhmtt/yrkstVFSJhte/+5Z0G133ld3/acV
KiYPIABnzM4OiygvK8EhNUZeCTcWOh8gcV48hBKKAI3WD5/vkbZZCEA14LCaDlaEaeHA6ae/3XEG
xAnDEgvhHPexCX4TpxLICeLazKOMzRZlK7pOCrkumOITzK+/V+Mh4twsRtJTHIg2MlJflADnmg9k
BZe8Z3G9eSU8Y/8En4kklV/crYyDToD6MFUaWHsfwJf4KcsjN2dIfGdBzRcwEHs+B0IvcEJTXTwh
yhZZ4ZoGIB/JR3oGRbdp/3LLhMbwI6/CywP6KpGRWCBUOQ3AhcR/god4uCaolSia6L2jxLQ5lLNT
IPO5sDQtv7Swx4yJYxGK8XVBIfzphkyOwDsnY6Zvn+cR64iZ58QuwRXkTOYdeXQ5KIXRdgwJgYRx
QdL1SqSdwNvPQXdWAWwBjV0nThxbgWGeWnUvscxNkUl4UCQKcEpynETbJ7+WTQ9g0U1Ixbw8CdEc
2UUUBoGNHUjuSF2JEAh2M03iSBWfk0dHuT3cVlrT7Ro4CpFxroNs/KUVFo28m6XLiEguTy7GxN7Y
PxO/5IHg3v2UIY4QVIzVLqmXc6zIU48N2c4Jq8jriCy/1iMl8JAJU54t0cMa8RY2GkncwiPwP/y/
6cv9GA3yhrN4oohkv90bGjqysU5YVdvEbR2ANKcUTo6IusldkBbo9pmq0OyXplgZ1zzUgBNcxXuf
5+NbijOrjgF3A9n1gJmn458mW/2dIEmvaCHLU5AxUid6d9S1B2sB0BNJ0fweAPxrLvV9JXoLQzJy
ED8f9ayP7h2kxkUd5CJYtwaVpWiNpS3vPutdQ17QCglrWQScxkNyEIWxSgGJMlM+p+PejQAXAG3A
wS43r5E0u/22hBl+ALuegdphX4RaY2c/gqe14njefS1IJPcT6wSNJw8j6yFnxf32ixm+4poLar4d
BMwflNDGGemuumO5vBW07nUSfhjADpuF3OsCJRdTTku4VhpQ4qSX1nqXnmE5qYGCztooLI6Em1rb
Ujvf+w/kcDiBnemGxUrfsJovsQPjWIWV4yDxvKw8jygKzhPIK2q60D3Bp5/7lt2xFHTSFK9WPyTj
GRfYt7jcNccjUCwMTTVCItvR5vJp9Ywrs3+SvgKSbW1KzOBGbH1oJfYRGG98ZQc+hsby8oQ9dCuJ
EYOUyohrKgs7FgKLhiUOEd+JA19LrT8pqSUe4kTaWU7M6uhAfrDVbMPrxSCO3yDmLbPE3BOoc8I5
tEiO0TWIL6oNH+1vNJiDGtla9SlYsaETGWyS7ZDq/Avw5K1IpJwOZE/9/mVyC9asDpCDPVswz8d0
VjpGz918qKF5IMyMg5N6NANKVWqy3T/NkBUOyo+uBkUJe1r5BJbu7nrg3vxvfFBjWjZc3s/hjzTb
w/YxPapp9rgRMNzFQbe4KzpVt6f1igPugDw7llL1H936i2fhVd5NLY2FuQGbVftKlrkLYjoOSf+a
o2xpJ4aFdBJpBE6dIB3lQ7ayeKEzuYgZbaE7s3nGbhUk9vB2P8VFovLMStov0nE1qxK5p0tOa5MI
9Lqrb+McnAINite/Iq0wyUpIFKRf7Cr9IWpYRyxawKgLhkENOxVRPIo6Uga2sgPRVHKYCPLqENOx
HdeLtMeEzUTuOR7Mx1bt0EUhsKwtjiHISZmYkRdOuOLq7q6iCk4/FevtA+zdrtREvGILNWPDR6EX
dlaqKV/EqzCYaTsbM6m2XAgK8YmSv2pmqRPb86DEz7rQkMBWOyt4whS0U9PXPXXLzwvBm5TYA3o8
x78RzpzOIh8wgBHyYPFFSKal23JvyD0ACjOJ1/l+9UbIC30aQuxiBpSUERu/hVWwKKAe8vKS52tT
uVWOi2Pj9PqugYvbAMyF5VT/OJpLuAMcAKc4Y7oN10emcp71cehLLaGXibnop3ZxivL6vj5IyYOX
Fk1M8HIOC1TkN9Kb9ei0PIQHQ43Q9uSPLYsBjI1m6Qm3PpnztIo/FQZ6dd0IqQijDrf/TCG2Amt1
IPkYt692aEqrosmZVdAgQgHdhdv/AEzTdq7vWdb14bQ8qMywYpgk3aCaOkAAkgrMzPfWtG1aFgJs
9KsCL/WsCl3y0eOfEM4yif3htbMxAtz0fimsOAI2+DP2WJRKQu7J5ttb1HWEoBsvIKMBaFFV1vIQ
Oj2BejdnMFs9Z3rkOqt040i7NN7Y3vJ5bodurcrpAYVXZdtdEEhyqdG06j5WGw8dytNEpXw7N0/E
rzUnusiDgP3OuVIZ+9U+CIAVzjH5Ahvi4D5b1IulghOQmn0v0gZ5aMXwA77xI7tJwLw/TH+1iiFG
qnI9Auojk5AAZVbTIXC4z8A4FK0Uvu6qZ8zwS7kEueOK/FhDGXNA3Y505lo63TzXbAZHy5kNm0YU
htENSAams+hklRaOX2D51sIHuRIpQvvvQOms3HRQ9+v5wCsZyIChkDSViLMlW40sDobUyPh1wCoj
BbP9hIty23VAnFogXSR7HTNO1eC+MkBV04w2PbJrLO/uF0gDx7yHnjIkKsYUTvQYVhZS2GQo4CEH
AaonTBca2Za2pTVdmysOtACSsEPqaT4D3PgfLiMzAcoFlTfKnSUqcLK9AOO8mQSUtvxIeX+TJuP0
PKqyj87810wFwhKIz+ItZj3V+O+qmOIHuFFn5D7kQ+7BP+97BzlGflHU9JN0zTQ9qoAN/I4xLImu
G7PADdqbTJwRv78X6UvhCaMnVN0Jis93iqU5+wMgnr9KDNZJo6ZhMc/SMO8watgpg0Urt+mkQm3I
OmgUrSOadnL4H8LgeUD3h4wj8+bYTYyE9teE5qCv7xdxjy7aihpbgqBVG8Tu7Y/SEXpNGM1p/C1S
VqB4vj2huANGdM6Z2JdudozrePOe29RGhVmRBAAsTzd4d2kyn5rss2XOvrQyYMz0O7MMWU0b84kc
Or8k5WoFzuoa+r/EUaxx8VFkTCG9HtYWMbN2fzPY15c+6dte/9yK+am1n9JD3btV35E20PD9hRLR
E6hLObwnLCUAKzR1PNfLsTJX0CR6Odil8bGutDZEAqDn7AK2qVvdSllcqN3nYbWHOfuXv1FJFx2U
sv226r/yHIugell8EeSJ3mN2K8mCN+hEgMzx4xZ5CAbWtGGwPOT3+iUW/dNJxdEuEezyz2NG7VfO
ZECZFYSGI3ZKagkaW6N2Q24U0rC4LhrMOHIaqYbXvZoH4Ku0YUYpbX7kyv59mM2w7vdmUV67zyZp
G+BPnAFWNO4AgGtkG2BAIEGam7FfUSCzXcnM8eHrTNGk8oJbjv6DvYX6UDD6HAvVkjBpmjluBptD
pOi7uwMYwLzgc0Dj17EGNmkzxp9oElqAhstEUO5JoBE+aXZXE09bYCJ7vhUwBpl9XbaKzZ8Xxv3f
u7vk+y/ou5meHUhdMeDmr4cX/r3TFL+8ZXhi0W/8PLbkqTtqYHrQGKLv04slwSRIaFpt29oXrEWU
psbmJFM1x1U+vaICK5eEX0k71QJqxM1FL98vW5zRxWQyjSrFd1r0Jqrk9ZShFWAjPJN0CVgMmkTV
clUZEbQacvXMucB8m9wVK6TBIyIHYeBJiV4078OgrT5+MVROMJ30ihGvfFvdwK2VXM2rqZ+JF//w
ep+0Al1gG9eb5utgvNkwj4PkuDwlgh6/lXxxQ6b6Koru8SI6dIANa0GfvKL+Ks/XZ4EVJKpv5EVJ
vYblXKfOtwZXxbT+6wkuGQS2NdYWfe9vJVOeyZECk9RTKx5MjXgWbDqnJe3vrYCHKyUWVERwKX2a
MiDoT9gQRv7Sp2HVF1raJMiMCkjQvEjlpUagLzhMursa6IIpl4LqwGnyyDFFqhHzHPw2tOJ0WDzW
MpsULLrxabTE0fWwK9B9Ej8Sk2q48aajiCvs5xv5HFAPC7xlpwXokyZYh3ZE8dtOefEFStD258qc
F7wJkYlbO16B89PF3OWsn5JD8wJKF9lA9q9xEjtOe7vXwrkgZESqxxQzN7Q84K51VaA/iwH7p244
RzGbvhzbHYkzVXqxFmMT8uoCXU6YObpsw6tcvF0zDRHNUNwM4tEEh1k3tSgspUyx+jZUJY3IfhPN
6NFdebXKFuB00DS6LR7hJyWqIBgHBmiIz+izuZjFgygYJlpOx4b6GqhVk1T+ToceSo27HeVrS4Q2
u+Qz2yi+g4zk7kz5mq4RbScHLU0/Voo3DnW4Exg9a9lOEbpxT899ngpiXINmsmEKa25Se7WQNkha
wUTsGV2ZwPmRiFh2TOB8wdA1VaqncmJO/RiQBcdokS/RWO+lzopttin9c4aZABdXCW5lib9yMZt5
XULJBCdqChYBjMS3fyGUK/WcSeiCLD6I8BrhYGq2GLznW9XQtjzbj6Q9nu2mzZRM6b7/Kz5rDtW1
SIbMPLK7JlSz/4cjupHbYttBlrsswPhGz+TyRJhrxaeZkrYh2JLTbM7KMd2pzkV3tjLwXUP+6s9s
GKllTpx5W51AsK0f06+COE7klJnWAzZUSdUKjqkBZg7QCizibLwErpmEDnuv80JCCGs9AhPK6OqU
xYNadlMUIHVo0zH2ezUCx8oWIEwYkvWeHHK6spJvlGcB/W6b6/diTibWltk/VJkz5zT3Oje/i+IP
vvtKsuiOLLh+m91lrF91zhTfwmeAQvLeA1Ja9cdyZ7gdUhFqz3BEcXhl+h7YwTTQIvCfPAlkMZDR
bqqKj6v27WXf1cI9ce3+NT2+fdhN2KXoTBURfpgoZ47X4rIq2pcWOT389sBSQZwOu8Sdic2IGWds
STzuktlRwKFDyX2VFvYCRmKgkRVBXocDffUcIWWPPbi3pbu4sA+H+U0bAJD/D6SICLLqeXM+sUj2
sX9qvKcdzaF4IVz6OPkuBOSLA6r68utEIVBGbFWdN9eSbTbzA5pUduxH+IOZyeDFQNHoyXk9zFPL
fUiZzxiJUCQaBs/RR7bSoHq0gk7OI6A0Rv4MDuC6AVdGW2dy12VIBmSl5ZXJ2xN0+6Y6CFmZwLJn
aCxICur8hFlbqgO7N4Lie/YSUZMSy+L8Ct7GxIvsttDjlCjXMS3mg5PT/3c1eHM5Ofb3oMLEsFu/
xD+csRmP0E2KsVVdmZwZalpJkH+8xVPChuclSs4y/OvpUTnf6WE5MLZ2gpMM2Nkr/poVHhHX8B+a
hIf3QGgiBSEtfaIoQybBq0kt0Sg9CIoOFyrR//rH5ctOkYFBrExeplXdzXdFjwXMd3fLS0VH0gn+
x6SAgULHYqWRFiM5h/IDh//ktlbx7537rnDXK3I7Rpb32xpXC2bNU3s+ItPCfm6S6M76ZwGy4cEm
u7R8RYl92d+naoRqKGd173kp6IBH14JUiEHNHTKNcMDkoDKuetXnnuRr0XaoYobr8RHssCg2nX9I
+ink/hpxWZb3VvLno4+VJNYebV/4wvwkNiDilPAX4aywBzLUZRdX+kOtpSUS+suC1MNoTT9IaOJA
nnJJgJGniLi8ZGa9TAEqzFjyBf5fw0glmM+mi39N1oND7KRdpIU0wRRcIspXHwkFrg+IUFBuGSvd
BGFnZ1weS/Hyx7gM+jBjS1yFMwPp8eVXFahEU8Y0lZpJv5TZubG/lsvoKOeqQnVfq0hCeIS9KPT3
f/Wn3NfwizsbVbYOFIQmu14UPYGW8Xjhm/rmjI6hxGK4keH9RO2uUw70RNupF+BdI+CkqGtFtHpD
DWn2sIDfEejNNNBIwpth5m9we8VJCegzWAbHpl7xJ5BjUpXVmVW/OG+Af23JjM6vQmEyZ0HHxI2v
qbrcfiCnBtcgb+riGydrJLu8FYrmPXFiteiTZQyDS++xMnwguHaGFvXso6OVhRUTH0zmAKpV2XJX
vWumvlUhUq1ZHkWB8DMykLDH2m6qPajm/Hk9qQJKMAbByyVAFqSA/B8hOS+XT485eir2WmPkNJzG
FhBJ3Nn7dj/vhIxUDCoh7KJau4DoN9Ke0b9mwHZFXsfYmBfoobt1SeT4+4+r/v3uGeuK4+Hd4Pyu
pdOe6lXTHKbQth4vkwua05SnmbZuN/omQux3OK5lYd9t80Y+FEOBFrMqvVk4zqr2V4DjM/Det7nR
APh2SzyjxoWmFKXc1Clen+eLGoHd5AFwl6MunWAwVcJEoRcw//6htfHBG1hJqJL+EmftdyoFqKnM
jG4T9tXGzPQbBY1Jrot2o0Sy5IxE0citH06dHqsIvBI2NJG7ZKsmN5s9FEN664mHUjPc0WhQ90f4
NBBaTYy98GMyoUSmc92HZYDGHQvBvVRq83gUvuTi5njHezWgqJcVk17vFymUfaSclFnZvkWv0YzL
1kMuCZA8y9fcIZi5R3ms0TbwA+5+iiv7UUMPLcS2tvsWcNV7MO28SNnqc5/7Ar9PKRijbr6wb6Zz
8obQeQLx1t427ly1OTfQry9g/gVm9MgJHnIOR+aT+D9/+qTk+6NEptvlu7pB23hjrYVs6uJysAWx
z4hvjigT3Sw/CmiArhDKsVECRAVKYu4S6U9TLXpFUsC7G3H5lFaeUYW8k73l/s3MZPO1LEf5rPLo
8aOnGkOZqeFgN0tjqInn3oxs8oeRLx+7riEYjusqckbDLjHKhWoS/gRX3cRMqV3wBlgC2pNNscxb
gjV8O4Ifdkya7CFB4Cgv0FkZTppEUjf7ca2jmPUWrkwspKA6ONbuA3+fz4P36IZ6CDJw3mjlEdEG
VCZP/+kD61CRkb4boIvnNLbndMZjQ9e3FsAus8on2EMDF6cAvFbIxJXuzCYhrQu98Gv6qZf7CwzZ
8KKFJXkSBszA/6v0wfeKUCWOWKHxyPFHR1AiFkvyFXaXzr5VxZeD+6zlNPf9GY1QUMAqEd2rd1I6
+wbHnkz7Qk9ZXS973ppRxNGldPmDvjo6GkqwI3kvixVsD5vP8cxl3poyVgW2LM49y9M98JGTwbmr
bI/la/oVgunVtF3KsiPGL3nj+XuBzm7+wEyQBBh6gbT1YlJADiX6Bcq6ZyZ31N9LkAb6fEHegibb
XLRI1qBs04w9M5uKgdXhkxDyYdqjUzQJi7JIn7XCYBxyaJn1NoJgOhWkjZFNzjlsYeWjWjZ0qlnt
6I4Dk6ZdSpBCNEkKtGHAG0bRNcYkWeBha4iCbBZhJc1+yyZ93V3Un8n7WapK80NfvbJPD5cbCHu4
D8S/dlwKEgeyYtqJ2im4KlCdoq3GRgqVNFC6yWDf0k+UImpthQPGEu5vt/Jina2KOCUYZxa7uDwL
mBDBjFgM9XzB3gUNtr0y12qu2jqn6Eb5VYJs08Qb42cCPmvweeIZlsb/EICTRHiq0Y1IUxiaYo/0
4xUJwwtAavpZBN24GkxvB1wAT4z/y/EetuydiRjuCjZmhlXBPBpKVrwidvhiDWFCS5fbftNfj5Sq
jdid4SQcg9ClM1HVbYb+n+lHPu1xr1D8dkp8clIb09+Sp92i6a8Xm9zSq/mdFkn8X/gVx47WV1aY
9miazC2swtqtH4C3ApAOKRwDa1E77C1oYmeS8jnTOgqmdLcuo8O5aroRjrKD6xv8MLkMStrAGKx8
adVl2Ow28YP9El70ciFQ/JPjgqrU2EN8okConBxiuRWtfxL5dxKOQ9fpUTJXX/mj5acTWEHZ0wax
4l+eMcEFwirBtUwEG8ZihJfR5ZI7/b2m3k6YomYe9OG05+xygndcBd7EbyOq6p8/uUaegIvCxIm2
/QZAFzoNKaADQ7ul44tIfSmIBIn6Nk3YhOcKKTh1xU892eyCjT8sZAX3s35n2RrePTtR5Qx5kagm
1kNWJv01NfL1w8U/yLi14vB5nEkhtg14uYeGtiwrzbZe/Na03sC59pcxR+hSbkz9h9lKE/gttOHg
8Nfgc1pj2l1joydryoLZvCUgKry0LvQE7g8Cf8tQWCZe1ntGfcs8DC5BKmm6jDi2NVdvmROWClmf
r8lV8S6vRJREboGYQERR6xJbQBpectss/Qp+nKN07nF3CSQgbDKJbwRGTEMlpqjfkrdrnfSHW0E4
vhPT1xrjsu8WDlcs720RU00Sy2zPnmgNw8PyNVTHR1KCVqlyOgz92HZCr0mHbXDHstjMy6k/YT3l
6FtA3OvAr+W886IlR2eChAtMhSE1mHHGxiefROQ14Wx8uxzS5M/73tCcTG5c1FiVA9ZZ09GChdIB
NEaduNSz10e7ThnGZ3vzI691UnM/VWl9iIJLftJBm3wgPxMy9hJ8BNQUJnggHIcRrLlVwF266m0w
Mmyq20C2SuSHGIXkmtTu1PHwupA+k/sBcI7DdC1lUvbwNOaA2G0WYT39QLxVVAN2w8bW3vR7FWKd
N5sOGwA+5kuptYULrOe+iVOdhFnbi5D7/fl1sPEFFz0LIyUNbWDKnmHLCnGAiGxjV3c4+VVODdM6
id6d17OJ8jgwzo5CuMW/Zj3POjfUssRBK0UlbFXdlLBZx1KAz1G+RJoxJ/0TbzWsWeI+zy8qVIC6
Js4Ds4Kq9WBlkuuNErX8Q+hUStRHE3i99v/urZLhiwg5UFAYnb6zSiRXs+FQ13Rmf0fd1WH4ukSJ
+yYm5AlP4ToIAgbv8c1fwyjBgwNPaxGDiV+jBgsPaCUphznnrh9jzCf5fF7xz3CXaeNyt04okCmT
mtGqqByb8lMvCmNagFJdqpQkO6WqX/pR0tSvnZII5BdgtE1S6/pTR6w7tf3yVno7bQunR+R4s7s0
LE1/uPTLqufsr3VDh7pGm18MRTN45nGNgMfPe2KwPD2z4hNNFfdjCHsygXX1+bq3gWCnnBru+WlU
JhQ1dtz95Of9n5Y0P/4cJwJ9FwmTo6S0H3HCX88M1v+iwuuyLuBYWL8uXereJpxyLWJhXHfSdiiO
t4yq7dE1P1rJaVpuHZe2ZXobakfiIDfROJenJZehQP2B6aGoAzIBgz56YM/nclxiAWWdrD1U2pmw
b/8FK41gWllEE/JMc+yYfqDpofDImb+Fki7MfsDxKpttwmcrke3j6je4cwTNPLQ7f4TH2WC93phJ
Eo9CTv3/2ZXh5esHZ5xVaRboFmWIEhRxFTQ655XyI3MJmnjha+awaO40I/n3QSwKTvC6rqkgK9e4
yeWkjdQL019eqxG8122ItgVnR8eMhyelutTnvE9OxxubInQYcEoofSlxouQGpNnxeISElpEx/E2o
YSX2M5T9lVt+DmK3Jt0HQEeQ7JIjx+7TWBvgD26MJ4O9RopiO6LrSQJRS2hlidunSlb8CsxJIqCm
S8MNk5y2rmjU+pqFFM0Sv9POct4/NC0hsHwkA9xr/35/9sbetRXFLR7rDYhFYEeYsbKA5fz7J9Lj
XTkJCVCGP9p9bwl8DplP9fLYneClkOt5k+JasTwYws4CMhb7OSoKsKuyUsNVc/Ev1GaLrjDcuZ+E
WwGZBo/c2YUeUNsCO2u7d0q+w8+LlgHiXjnyg7zB5F1TyPslhJl6jzrEmlU3gLxWrrvPE1EpAUo+
AcFBILbbysDdw3czxOVCGMRmLS8frH7+lHz7tbWj4V9Vvf5b5iN1OKQ2gc0RK81Ia70jxej53Wl8
FxKm5/0VmFjHg17cIT5BO1kPOlAYH/xLmwSq11SK9d0q0VkRWhb1i6I+MParwVdBhO6PxfxuvoQ/
36JSKzBiqKADDqzCHaBtJkCGqYFzG2Ez7zNjic8yyDFHSk8g1bFxsBKlv3DCdW2FpNLeRXxeAPsF
CMTobu49a2XnWSzCED32eG2QEBEgRpOvs59gvKfvMIgCzZxRZnwi8mFClJQXkcG3s4pWbJjeKpJz
vBq7sKHKmCnU060ZDgtyFFc/vdfeLIZPyvPr8HVGBvqdV0HNCJXYx6zd5ty7bxkOMAFzPoHGCaGu
N2K2cmahmGU720Ey++n99Mooo9kvqMT9zyXVYjNfN+SbWSDQPeKbP13zaFkH1AqIKNt3aX7gGUdd
I2kXVntGJ3vdnMlJ03ZcZNlHk9DdsR5LZ2m4awr6EC40Lr9V2r+L3uS8MjlXwWp8wFSGrPGwJ5um
0ln3Vnhf9vMz19gTKDhFSnif4e6zm0477mlKI9okt+ePFvicUZJluLWh1nODSNUESkgu3uRlzf1Q
ZWwLYkBpDPqGkkiBnme27Mz+NvrpUvUUT2x1vzXZCZW824FpS5A+3WNJUOOMMvxhQEQXc2M5mjUq
VShlQwqTssPr6KntdU8UAkdkEVthed34eIyMZQkE//C9Ap1m9wuooCe1xs2O/ObGo6nOf8vRJQJ4
ZC17gg9P2xdR94NoMR7AFlweYZTC4yjX1SA1L05v3vjhBYQMY9VH8AAgsDI2EEP4fXG4L5VGztBe
rM9yrzqyiCb77UmQcgONUpEHr6B9PteBRX/1+hoGROC1ddfxpeQS0aNaDTSS72raRymmi0Q/5px0
bzhvesON1GeX9DVsOuf4p+GlxyWyfNu8IaSLJDfAnw4MKoH+Wvyvq0iGvH/sPbBZI9oUBkpl5+68
8tZfHPYb3jubRq0hGcTjvzFf4MyPtLf+0m/2bc1a0UU5ibfeQ9kL+sBeH6rheX0WXo56DzOZJGkh
xYzuqyi/dv46NNksZPwTPNYHc0KSoVxTo344N2fbfJ8WNtesnOhrIhs4K2cxbxRVjN8Zv2mMMfsg
NB+9xBXOW9UNZlZH5zQ8vHI+b5XhCm3kqcZJhEHWB+2ax/LpL0xdJrxYsTMVAKM22o8pseyWHldc
9+2Bqq1uh/jEV4bzU0S+cWff1Y4GKr5Ehzjbu1Pbma7YBHH2J7Fxl2Uz+FjBxiFpPbn6LzpmO1gT
mCBpJFNetXelb0CM+XCQHbvduHW83L6ra53rJCug2p9tCp2bLUBkWVfqMNFCCxeJzWqC4MaI7N9B
2cMM+yQ8w4sdjCSBd3Skta4AtJJmhkL5b4mKB1HNaL3QP3IgdJaHX7127k2RALV3VYg8RkpJ7Qep
/TLxi/9hLBBcXtRYA4DIOpDOGU4B0zMZCiv71DWUFjyldoCuQN9BBTYDpoWgY4rdYq5zN3jfl71P
3fCtLjqlQBQFvIQEWcd1kh6qG9ygzJmLWn7vcoB9z7q5lwqquDd7zDme3pYgKNIu8/azjKG75lFn
4G3vVKQJsKOMh4G8y9bXwoIKNlvxIHiec75iKKn24aBMuwnMh1O9PEEl6DNvka8JjkAVjE6qoSkZ
sPs2+KMFfQTzo7XMNB29e80DzX/9igaJf39qLTZsfczFp+Xf//R+VD5VUWxv7HCDhFVIudlTWhke
lpwJURZWdK94bJe+IHyYeJlI9aXj+k34t1B1pU81WicX6f8bafhfW+ThRtJWVadmN8sJWIO033P2
LQq2QgnbdL/icUoDDxMFilQFBPcFcaXo9Yj3xV2FyhlJPIiHEW9OyTMtlTqtLLsX+lkc3ivY09FF
IiGQ9bYRhtcN0nPSzgLDoPBMzHDKrguk288ibjFJI+EanDaC85zrP87W3x7paEWqFjUbb/R5CM0W
CWpk1pVT8GqjrtjngxsOczPT3OGC7+uIG2NO3E//XV5yCShaI8tq40jIVXad/4uAEHUzUzRt2IcD
sjni+BqX3CgODVMaoRnzp0YuPR4eyX37DxpBR9gWFOPWyBGM2Ax9eYhXIf7ZgcqKnSw/2mpqi8fd
BnN0RMZaB98ocodd+SYedW1qZ32haPriNbc3UpY2MbC/C01yqhRVmkrUc6iZ/F77oMcbnpTmcMVW
OpEtWnceLcoBQ3yg5ua2K28B5aF3Aq5Avcq8qPfjZXarMWs9drpPOsFhQfAtx50jTRKybcW2yzEd
1ZyFld3/KnqzF8z/E5092VKf/3KH84wJTJVomf7YMgGcIxds708FsTXw+UnHo+o4tg2zvlRocYlb
Ng0kBIDbO4DdEtBMWaBrkAIXgasYEguTPDRmfLNxqQxurhNzTSTAORmPtL8QV5ofmG4sOkFN4XEG
SKfMBQ10+DzUhmIYtLo56IPCPS4ILd6DPHG3ytprMo/B019tmDI6Go+WBJycNhagkkvPqsVe8FG8
IzHDOvctM5mbjb2omV7cSTefnEq3gOH3rGmagkAW7iu3mr551l7Hw60qziK1dIziJIGT7DeN2Bpp
ywJ+h7ypCOHNC9gD8/fhfRsVnlP5qDK4iZU33azibWp/7rXpkE90GkPpic6CUKf4McT3EHPlOJEi
byGFXRQJw7AtyYKX9HGWCBce7auquiwa2hpfkW4Ov4NhbpGhHJe+U+JL1ej0c4FgynottFFiuFYk
vqPPUBBg9yokIhfT2nFOG9Exg0zfkGOpxPG18jRQ+0poLVCGxH1A3rPFN/IUkQvR72xtGLjQr1Z+
sE1Ds8m3W8VsRXLTWSsLEV/zWilLIqqCoeTDDLnHa936WQdvpdSDTYxmiCduaj8elE6+3ekXC1kz
mc2r66MdHEalh4nn6Vgg57dOQC6WzlmFabijDGTLPsR1iDZEscSOl1lB7JXWoKlKd/XkDu4QO8V0
Y7hXqVuSIIjVKt+7zLg5TyD0f9o6z7flOkoZmc9S0NoBPpj3lvhvjHuAduwcFnTdoyrCy6rZ7c0T
mfvbf10U78X/GK8QufpeejGpihF4ZGBDlfZTps1w+6FEHZ7XckpnJXNcL/XvgYy9UTQbibFbgSj4
JSOBcrEj64JuVGC+N4nv3zaN/FssaBQywwUKOFw1ku/5qlUJN81fl6t8R9ZP+cYeFnHVSWFIdB2S
NafGxkF6KmIO154JYQfWqdLMW8uYUp1YFYK/lrmLtYRRxKEB7+jEd2eakUesB4LtiujswK4l+O1A
DQLsav/x0bCdnlzQZtdj4cAbJupyELpDMqe/35GhkYTiorwtIFeLc+ik63MWSTSdH/8jqz//z/cK
K31d++EjkNQQci0YO8wm5jL51c7ETFLasU97QjQUFLY6x1KTaB+zh5468qU9wuqZ+uE9m9iEz9QQ
ln46ZflZzGs8928D3ECihG8uD3mLJoNhQUEtiGXm6/IWzDU8EuQmCpjpD2SMao46q3be2zeEvT7w
arYD7C/rqkk6iAa2Szc4rDspBbxZqhkojdtXOpmGnNUmqeTKXv+Qxize8d8eiE/lzfVhcKHIK80V
PW257Rp7Oc2bo0GiiFIRn2dok9GuNKtZNZxa4bUlIaSPCUmg/trHClGwZpDywND4txpfhuoTsUG8
5Mfogypluf8HwumDeOnqW28BB7t0fIeOjkpRePef0S0N5sa5ngJs4os09fO8XqZ7xBF33PupUZWK
HoC//MUYDn3U4lCODgOALc3ZYFVFHcsFTo1IaCrGRetYRqOwZa2Sfb2Tu7X/J17EhIni6HUqx87v
MWsNTb/zS/f4hPx9MeOMjczYCMtqJ+X8JT8VBV5ci4Gxvb54i4wzpFF1TqFqAzPjyiOgS22CbSFY
J2XxdbAv8KKVrF2elpq/8MkyWmMGI64fbMSonvD0vCBsbjsaygPsdADsBs32tWQitBe83iK3IKTw
8OFfBGyWR5FRGabyAjtKw9DbCQNOtZX0hYADY6nSmhm6YGFFuvS0AY5SjQV02/0MN7tEGlGANy2e
2XaLrUgcLyw3iwzJsByCuQaHMQk+ZkKc6j22fvC7lyhCY4YW3zvTbGQPBfgTkKifq6JUp8o/nY65
RSbwor3cq4dQw+QZlZz6PXZytEaM2CCsw3dDDUbzxD8tEHBh0UUNHwhgx+tz0Q5Uf0mkLiyRKZx5
nlUIvJeH8J8FQTLCV6ETVEixuiuire4Iw1kuGf5fvoCn5gUptaG8nN9EzpLoWVSxLBNCoxP1Potb
oTExiKngOj4z73Z/JAH82SqYDABwM7cmIyW+Sw/+PuaGoZT+Zwq+F6cdMI7dYnSr2ZEavt7TmIRw
p6gGG0+O1ZTzVVatkLInBs4DQBBWe7E2QvR44z9QtHS6rO+N+NxWuKOV2BoDsySwxrDANScIWR40
VhglUTB+W4bmQAL3rPsVnWlbLIHwhFvFRX1nhX01AtySjWeWXxUb21aRFpGk0t6KGiU1bjAotBpu
wjG6hlq2VO9v2kBZfYzRph43Ay2IPcA+Y7phWXOBQCorrIcFmKw7AWdwiCbyLKPtsj/Jq45Czpgi
/B1EtBKM7FiMHKWQrNJ0TDCT63wEQLwCSYp2cOqjNVzjYsF2vsXTq4F/q/835MV9+KUKNwrCBSWc
MzUQ8VXSn9Ua70op7fUnaBJ2dRQ4NwhepUeaBhfwvFrtCE0FqNIy7lvA2JDpyRzAHYmXTREoj5qR
mFSLvn/bZgus1KQ8nLfAbkKpFV4rkGuLM1H8SAT4Yz4I26Dt5qitkq+pXFjgEi+fHweZg5sD19/J
PWUWkRm7A8RJCas5NqolF7NK1Wk6B4z4dN2Aaa3yGMOEGUPs8AsOGZ2Azq2SCptSzvOvQaAp4YWd
Ob31BjTXkUfKZ7ioz1kEJg5jSNHPgllqIqUBhtHsGA7yXxJbCDMrFwpyl6KWPwcuTahnczxV2Ayu
1swcF7+q4COcKZJpRnSg7EG7iOQD5ERR5GMKar02/Oq/+/Jn4XIuWWLnpmUANcnhYO5oRCqcW63/
yMOOn5hje+oID3VD3ayLjQnSS3/jgLGC3hiIQXPlHXxcQGnUyKTAxXgxB/4BarRH5/UCAOPftnwc
OCw2GOxJSPsSKsjAXHH0KYvk7IeMpTwqXex2O7ESbVyeqUKpEBJ4XFdp60vL/sS7du8XmTKHqq28
ZR/4E/ho4cfgIEomUc80f4KjM6Kd2ELADnpZ1M8s3yIemoyZ7A5F3ltn6BKEsa9d0yi0czN5DpzB
fIN/D3+eRGYN+SBbU+DHhcpXQx8Kc8ZenDeJVzCtYxgc3JyR9H1oelt7M3MOyChVuI1UXujS7wR8
nynaNs4hbjtk5JrlKi+bmtyKF2JOR3VlsUj2kssNZ0uHn9L/npZcHOLR40ElH+p5IY/z/BNYiWrs
oLxN0tlZdyypIPO496sffQoUPG8VBKE0A3m0xd8MVsu2thXWP5YtLIgcLKxSf+xoTBKVrCpahgBw
00BtpftXwSY8M/rQJPZ+zRbcscHCof/qX63Rg342QubTMo7FjXZnSN7fpPbrFvnidCnAq4tAY0g0
gqgELo3ScrukQisM39ouZA2fvBprT0EkjmtWxBTXaWalJUmMGKrHBUQUGIoQC6tIKA712v6jhEUJ
dFcx65ueVro5YolegNgWob2VIfnl9rC4I7b8sAo51sPSN6f0L9r5RJ6qlbno+QjU8ZnxnVsnxIfc
Xfvt3MvQMfF0KWT+B0YDXsphTTSFLN3dK58oFPzeorjBuu6svBr0rFyIAi24fOV4/FmkuollDTwC
TGE79fNBQmcP1XOKO7y0J3Warf4YuN2HIMYmmiNCHKB2s1XR8gJKtcFm4URe2we3QsNzt48v9uoU
WQKc3Eej/Prm1zMzsrCgrS9F1yfTi9B8fk8z1HflvF9k9dOuTqotKqlAeDwk1bfH8lmcKLMnV0nU
Y/iX4IgfBcapzdQbcCr33DMgYqhgoYkvW2p4xynDCNsYtKPWFsooms4WcWQgMh1DnKpGIIHLMg9G
UJOnZhMSVdcsPHq6cZxnexvS2T4qxW7vLmuYb6Qjd0IWEpkxfXjHqreziR7kIGvG1AmUscl6gk4R
qyBAPKMTdA0SRJz37teT8gnfOPuL7HL/P+uw2Vkr1RB31lrDEb+On+sThZFcAWikZBqUKl8WmaVu
Z8CxFqLLxdnSCNUX0zwialLxTIIdTNa47uolA7xg53eWQ6xTFKHKLrptLbstzFX0/QsdQH831uWG
O4iM2TGyPbkll+x63kv2x4FkFIliTNH87dYVaO0SMlhjX++mj+SzdLZ5QvDsnfi9Mpyvex2ybBtd
huNCKc+O2W/GsjFiBQzr+64Q9z+kx2E2+A4X//UV17Afl2hgOjgQE1VODwvsVS6e69CGs091ZKrb
6XnOqFDIGv0zpdEGkKTf5fUcsl1mYYo99J8iXM6wwJmKbEcJhhj09FuM24vZBcL3R46BBPCTVXCL
xka5VtePjr238h/zEHZn5h8MVqU6yACK9ek4G8HZZg/xuFOklOF7o+hNa9kh2EprrdlwCTaG0ffR
Gay5XChmvpnSP0FcR8IHKe8MH5D+RaWJfzqOyvOb7j1muica4Ne7lN3v8cMc6myx4FX1mrElZiPt
IQD+pVJ5Pn2Ub688NQSqo/MdX3al2FQbqDspTvdnoQJ79fyhFZKI7k68BnWmDe+0QADWn8EiD5KE
stoQ8PamXTZO7zovgbEbrFCbnjcQuRysfb8PLhpAMtefe6OHK4c+ZbTyG31m0JUoILRsxTxihBHA
j2KTJ9lvkXpRW8O/lfFEWzNMPD1ZlU28731qQJ/9SFZtMXfoSx8UB03A+TPxbt9K76+SjjK1V6ku
kmruPXYHVSklgNlNbFbySN0WUyEmkSJauq8lFcLzkvQpRJv8JzMCDnNzZzm6hvF5e2TldtDy2+A0
z+iYFjSUbcp6eswLefU5QtZeQibpHr0s13HyZnCagUJTI+t7j19ewsbLIY48Zxy55kPFwlQF86dp
s4fBLqx1+gqn/XUISzXX1kPFZTuht+kx8DWZZQNwzaCPfQuDCzEkGH3p+ao8oC3e2zS2ngFL8eUL
gopiJLKzeQPb77j2bvPsrZKfuf/PYNS3HeeaIMB9oAxe+723NXcZ3CFcFvYexONoPDqvOQVcoq1Z
V6sj7QVauUH9gl3W0wDm+sAiWuzwsezCKss6xeQWcZ972G1imIylGU8Kgo6hhMAo8/i/Qay2EtfE
XuXDngYSwbhzz1YKT45KIXN/tL3veOoQg6NFE6BFjepfocEjsHQoB9vlCXjEsqgd5gru14XBziCt
yTVJB6n8e/Wf2YqCYkM0L4r5vPzv5qR0S6Kn9Kjej+i7ghg/3FVtqaJkrV9v9/UwtlcoHGJzec0g
Dd9SSmvL6RjNn+/gg9+P4gy+Va5L3n5qnM231ghlvLml1q8hC9ddFXDhArTwUMiuB1oIuPi5urRm
d3pRKjsUjIa6N36ahITfUmbsKRAX2qkHtsXMZSwb+d1PfI1771Cv9Xq9pWEpN+cmFpmZdAgvGdOm
7F0KgerPZCwFej7ZOkQ0JgDoL81kki7E1lqts40RrQmhzU3EZPbnp0/r5Q6s4YMXJFbkurcVYQmR
T6ZYcjl5Bn+HOhSIJOw16t418LRznZTQ7WRty+cAm8w7fk7ZnlaWHcZpQOe0B2V6WT4ORxWNMBcT
jl8U4JxYOhP/Jw1Yw2o9TGnkvEWMku6bl/GfYZpEFYD44Syf24SXkT8pzOEBWRlWe/HNCr2X8gIP
8Dfxcwp50xkrR7GD5Dc5xnPPx9dZY02UVQwuxyqHymP+Z688RB4zmsi+K8q3wOLCS2FDETNNnggL
M72PK0iHsbgOc5QoHzfHyVwHsUQKm1ayy1WA1cmNP3nWhG/8XxCmddKcN4USN9IuUWBckOEX6NA7
D4EX5PuJn4RlE6qLU5Tx0XGwfRBVIDWESwcbNh+TVsjafvzIfkC6v6jaVXuRb9eaNK2dsLhAMvS/
69nkVCSQhrjjnrFR5d61amL8bqBvpzWCm4Y4DL5EfgGtbqTQX+b+eTFqHORF1Nlzo3/AnNwJ79Ae
rEUFpsVU17ZC/gDqtKh3XKRwI+Koqlu0uohHNaNOeo0MYxLLbyijuM9n6AP5VYPd2OpRl2ThSBVz
IvooqmEXUOQTsw96W/puUjj7PlxjUNpX8TN4yavttqFrsn5E+Lwme5nUcqqX/rL6r3vSLnQL8JbN
W3Eh6N6s3zehzpnuI+u2jojpeiNuuSdKxDUYsaZRvjMzfH9McUX6x5ntQka5lN59fUWx1ByXcrMP
eizRGwuqSfqPK9c5DrpSlnwYxrBSaPOvtfihDz/CDMmgCva2oBpxN+LzJCNWEkBg3epPjbguqccN
gsBfEzsSe5WY/4y8xRobP0FgVV1a/k5R1Y0c5d34befzhK/zuy2/2OndOxkKKmOCtCF/XGegq/Fh
VuLNey/fKhV4eivRjKtO+arZRWi7q3q3NhAz3mzvGa1t1zWm+b7PLbYaqGBGjp1Q28V9d0PrO6sP
rsliPdxjfOoPltCpWj9ChyaMZe0QVZziRB1GUcBer82vHHywiSJqlYwrmrgKK8Vt1TrkS/JkvB+Z
PARkdIbLuB+gCS12Ed06jJ4b+3/85nD2gZRyyYG6Aao/XEi8aCRYNzw/CME8Ad2ju/cGUmACqste
ReqaR9Bz/6+Lm1d95dg2CUiVDrMxKyu66EZL7vdiAZhICXuLnvpvqlmt+aGhcXIJG/7pvnB+HbQ3
HA5GLr0ZCBsDuObJow2WndvMBcTPnYyi1gLgs4sJs7+gWStEnAHs02baUSd1l9PDBJWmjsUgnwNM
BIb90S+4fVCJevM4JYbcgaX4K4TLBrd2oiRP/QmESHZaxxIV4dVg747nrA6SPQlH61NCnwN6BV8R
LlGZlhhzWzA3wJ1i6nSG4THSak4Ff692oiq1uweVnis/T9vuN82mJ9JwjXmcYYrxBz9l+NAMFUAc
WXTR7TJS0cns4bkkqPQr+gC83SXmYGkoy6xY1V3WOVIyT1BYpeOXDDdXqshymlDsxOXl1y5+iMYW
GE+bQH7wy+URXdoFHrjV/B7ot0DPUtEjZ6C9KIfu85DVyM4aDyH+L9Ak7FB1hxsppXTZhLuwPFBz
FVlmR84Ad0n6McfOdHvprVk60xNTIIPG0GHkdIVJyy2mC7f1SamDPo0Do+02toI9FWN89NsanFoK
irbruMgNNlkhx97kookp7QFSsoHidXGulwK2ZAzHygC/wapauYQioijwlxpeXx9mn0W4nKL4HOWx
J2oTToUlHsC3R0mPscCbEKaReapfZ7WgJFmvyXrsRrc6+1pJMt7Dilo20ZCsNY8zwfK7Y0d01mkR
ZsWSv7/WwEVyAcg2lN+6jtEP2Rh/+wbcGcDy83tCoiJOGMHPJEBKhcukzTxEEIh1KzteTyCTobtC
Cu2VS8np85C/LxYAKmPh6T0nB3YKsepxL49x26wzc3XfMwzXJjA2mgkRcD5HebWv5z+7X712CmFW
KtxMW950gekFYPPJW7yUZUEfSArRL4DztYkcM6Zh8NFhRLjwYh+4wp2RGMco6A3dhWof6z0eRhCT
cEr6gI6+jRI+6yF0QfRsTDcSbwjBQunUsYcAXlEvZt/+VLQne5nUH9Ge2mKZA0bbj4qCYv0Mfuji
qe4/dCxLy74HgeP5jyIZZ4rQsA0KfliLfYOJlIeAnbzr3U4Q+6ysojkFlIcCx/UoHIjvwC9IEcHS
8ZPcEEjYPr3U8vSffffp3FizxVHI3S9CVabH8xApbImNEZ4d8Nmw71q5E6joSuEx/GfG4MWCeZgb
7rbPoLIrxEkk6FZ9z9Ehn/TCupWSduW6fOCh69J32qix/p/AOPbY12XBCwnGuT7b3P60nYUcj1KA
HiQMik+1lcwwIJpHZJGadsZoRuKTrSn+Ibz/Qrrqqy1QyEAF/W+5o5AnenVyE4yBwhMU7+m4soQe
a87lXu/8AlgftRZBLW1bddrx0bneHgMcBC6finuXNjXhQ7P1YxkVF+wiZ9xGZtCYovinlSE02+Hk
UC9xwuj2PygBUMI+L3Rdtmr/z9s/hsKHFFS2ZhM7sh20Cmlz/fHdzNeZcl7s+Dsx0f44u5adHrS5
3fwxFKQHozaQQBcm0PQPVi2yoH/lpJ2XNlcN2aqPkD0Aujn/gxQlECVaCWw2BcIYQUfGCm1fEkAc
ohUScBmW8StzKRNOIemsQtVMQNiQzbi21gL6Pkn9Y9sN/pcfmj59aXSXTHxLMQ9cxwwpN9AxayIE
fLlSF4Se81TuX474/KW7I+xDJV2NFlcwksdhWsBRicnPqC2/FPyz6tB0nzcSy1HK1B/4CD6Exrkj
Ai4Xqz0dPkckfJjyjfDHzAEph0L6KjoTxTZ02eCtt2PiGCj7qSsJCfx6ZCFtCDgI9KKzPmKhnoeb
LJSADOBSM5RIDnnyQKuzuZs8b/j1bSCbopDVwV471u/hJobCp74x6eDEZAR7GCsL0k3Te63nYD2z
lcqlw/y82R7NK2AAk8h0SUQkZ7oYUltX8ec4jMAEAOfwEkAwswOWPFCgIY7gZ1LKOm05AUeYBgB7
inloQIMbAPj19ah5zCTsK5sIc4HM4q8Ry0r2UWxHAIcjJcyPlL4A2y/6Ppp0imD+RXLxu4A2eKGx
C2YpqKfFuyKrOVsJftxQCABuK68SrVSQRUYXr906XhwKVIwwM2CXmzR8hS10nwHQKm6Pk48dvBrd
V8yPnoISY+nsCgiQ+F144zN06IjZFL/vReePwfBuyXdmKHYl1PILvepU0rVAXh7oIsMpJEM1at5g
OwuW1O7b1pfBq3vpk01EIXpJ4NYmCRnOBy54GWYxjnZzBNIScattwS3jP06p3I9E7BcspNlV55lp
hx/iE9XRRayFj0LxhpTxQhnDPQ02HFu+dWWpTCVMSEGbnPF8GHstWTjYwTX55dEl8hhU3jHAVeOp
+8EZsSUUnwjezqyMR/ECAU3Ber6k1lYGOYDZ0MaRgtnhGe2ihZ7cj8linCGDPyYLdRJnREv0akhl
Q0HBhEAt2Qdvwra3s+5GApiotskkNLmlG01IsCTTU8SvwgTsLY2NeYr/Xh956qXJcqfJa39FGDCI
pFRUN9bWS7kkk00K5ZBQNZstNLo9uRBh1N3XzCpSzPx1wO4ak/xEHlOMcT6qCpPvf5Tb90SyLfjv
cjuMACj5U95WOAnuGtXhg27GXckcCsCP3CF2cQ70TzLzDaKNU/Ws5P4mfbt7XDQ00YXQJY8+eH/g
+vjnObNAdgZo3JxuZVXanRPDLtbbdLqlQOF68jw2qMyYlQ/Ufp+WuS9iC7TKtvO1wXO644QDU0Gq
cwKmIUyh8QO7LEIO+QMid35r8dC6rlulXFPVuo4f01GAajTlOvTT6APD8mUf38Abu+pb6srZYzWj
v6vvbKV5MNa9Amdkjwt+EnT4jNx8hY5ZYp3FsZpfvU0gzBX7p0KabUCeoDzuNuoWrVFxOHPj3fGw
WQ01jX+nSx6lC0s3CzMqmj1ihmlDWx6pbHRHRakgbi/8UfhF/yMYbaAi6DKFUzwt9ktmvgUDIZ0r
5ZKPYivI6n4g205RtmENGvW4yQewQPAkExK+r7kwdVYMFFL2JL5iyiBq/pd0zGxJTiTzjn4NHGHo
vDpmOiz3qtI4a6hbPlXFRLnUtfzYIJv2og2RE9x2fbW69HlWEHnSI9+reuZP8FlBgKdSACQxcEHs
Rbn+kzE0DNhJ5lkdTLqVKN3mkvIlLANrJbla+EOmbHs7JCLk148Z2EnHs8BqlGPH8fM/Fw0pq6wT
UJiAYUHB7Rr2DbSDTk3X0d/4bYEXF9p7OHoFyVeBjxd4UA1lFC1JVBSJA/No/1z//9beG98j9gVw
fkxi5DO3tgBtqA23IhS6bobdSjXj1DqaLNeHqhA8/+AlObDzhgM4JRT1pEFW5RL3LdoZ2NTtHUOO
Wq7PH1S+3aRPN3IL8jhrwif2cPNoaY78G6tbMt7wZ+uk/ySjQm95EYYr5W3Lt3AHSB9bGjGmNQFR
PX3CFgZGd629Sur7Uqd/uO9YAWMc6Z4TcSqqyPK4KvbsAeBLHEoq+T+fgeEityWh/VTYoSx7Ewxe
edQoa6tonNbB3gxLx0iYqR2yJpAybc8BUdQNY1Jb/qFR3lZbOxHckucOzoMxD9P3gJmO7bBJf6dw
VHVvaYb80F5wdrO9Vw6GfwwbuQZJsNjtqOUCp9Lbi1xtddWhbEnkskoToeybit1S81RWldIvLo+O
IwYw3jO9oNSfTKfvgHJi06+cMa2iN7LKeU7Pru4bQ2jy3vT40bvdWyG3spSuX9FCcGIbb/NDUrI/
P1/FbwVgGI4/RRAquvqJkicGlIj0RDkxnRibTqLB73xTlfFhPo9LmdQyUh4T+OohagMsTxJHwLD3
8H10MDFmdMnQWcMrENgFM0xWzMz7JK1L4en/CLPF7jm05UgdF5bhJmcafI8tq76IfQnGPqDe9G5l
ePTQ422YwfYgbG0+0QJafqRsU9rk3HaB1gtEiDGd05LULZw4jxzF6aOR7q+gFvIUk5q750iJrfOf
29/p7rBywS1efZEH8e3umUhk4GfkYJ9VwdMpJWWaaKQxVsKGTvAYH8IaAaWNKzRbn25xh7kLf0RR
nl7yFo0KIMRmc70wHkKMe15z9Xe9dcBXljNsfmTNuQkrJXc3yaGOx3kbNRaTz1yN0EgxBN2HZus+
x1SnEvZFBSMQotUz4cPBK8LqorJuPdgLuR4thVa1XwjnKJA2jvcoyjvVdZfsM/G/WaRzFfsPyenM
Qjgh+MfpeMggldHx/hhPeSyYsi16oJ5mEaC0fWY3Y1EN5brDgnztODgfGL8DI+kgVZbch8hT1CBx
23V1ZYX4AznNd3Qg2MQKNBOTj7sn0+IKQmHFRlpr90KEZAhcYn0HrWuQnTye7Y6CwFe1ziWXsjjA
yx27uvVJXbh+XUt2GMQ32pCeVnB9J4dgdYXZd6w4rejtAIbVy1Lf+qel8t1Vs1a4tRIrff+QcHPz
2ItWiaNqLooLZjfzQe4hF0j2bt0VsQb7IWtiL7DDx7w0BoZfXDRoSBW0YLN0/kjNM/Rx31MmY0Q4
lbFvDqE0SJNBK7C80ld6+OU+/T3k6YNnUHtmEwZsPLdLVrmotg3Lt/iSbX8TWnvRmcL2hS+YQeg6
al+lvYO7dElNs4MNUVxdoghIwBJQo9FdEzr0HS5bGS7M4cYBXe/bM+M2lGza/GJK+oCu8dq4hg+2
OSuBT7o8q8l2e6BP4CTPeEM5CLpI7b4NygugDtnXP6PM/HhDek02ZG3+SKoXNL5RzfBD2i4zVpo/
Djlr5jjmyiYdPtA6keUz+2udpqdHsqyh2/e/8XxhM2zcuLR1jrWPPzWtcdF40zml+jur7RNw+cc6
XAk/VBhHKQ1IIcc21LjskXpQIdLprVQYTowCmY8QxGVQLw+7FJjZREt9UI5GTZWBUEI6A0nQ7Sp5
7eCRM1XYRl3MO9tg817R/SUqtwoWjyG8PgaR5p1B1bAL512X0rpliWg0B4fCVO1W3n+Ydww88Gxy
axJqC9/VVt84DyfPZ2UErJ++T1ZFo7SsK49WxY2Y5bnYDUfh6RhHuWEBd4X9JIAI2r4MIfHPsiZu
an249+idIhWNMF1mawVo+0/Z3VcDJsQcKeegwwNrEO+jKJnsrLWKSjp6i1Mo7/9VNMfFZsEQ5/PZ
X5BvNlhLizLrIzLapthG8U2VcZoqUKKlLkAsobPIiyniXbX5WmcYpWXev8VUi+OWlIHJM392aO8w
DrewJT2mzXqLnP3cCvg0rK3CZ2l04Ho0t68BRxC7bcikBGDXee/NW13NdbA/FeIE0ge2LErbEc6F
E9t9BEX8K4OqPoF3XeCbS6AIjWX9W40FKErnMqERa3MX7ggQeSppU/xLKmc1Do12H4SE1p9arABG
GMbVAr8NQ/hIrrHVBOlfBVFf6n+sLIEviqU1sTmtxbhYTgA9nyd6VtS3oJXoVoPoefOnMapZDBpl
snthqqpqEqQRhoelwL2H4dlR/O+uaWUnHbejnm5qZfnxxXZH0nfWn2PmFwt32baP9Pk8yUc89g34
IWYCXF67VjxyqVvFeE6Er8nsebTq2D+NJ2JGNEe0W6fE1aK6B6Or1BqAgsdHaQb9MxeKWGW732u7
HdnqAkM0SZQr2yrH02xljdck1ir1QShBlaJzXXhC7FZfeyZSI9HlQDa25/GIiDQmY4uF+rdfGiDh
Mvz+8HaGlzQSvbibLDyh1AsPisawItSYH1wwalHwYbqKFUSFqVGtQtmWDAoGhXCAKO8rgp2Ix99X
3YAdM/vjET2Bby0OSOmEWagEsc7kxnBwuOkaUyllgqmm/qr4lg3rL0/u9GejRYpAqFihnE+x+Uky
pMs8GjJIadXRiLh3l/Ke15p1WMYbaTUo8aR3pXAkrmkMEf6i5hKh0AHzjmC9UQmPQV4qfXTiPGML
BXhkETDYbROFtqlVFTh+UlB93emq8DCdpsJ6/K18cqFEaEgNB+67QjDHH8S2ywWQ4CuKlMBNYe/Z
PayffNaselD1OogCYz/U8u085Ywdc+LO6KYhysIoDM70w1qirpmW5I/BXK4dz0jffFFCgCxVHEee
WkYb9LxZq6Lhs+ISztUJK34T/Aj/fXt3xb8WDdicvj2vIkr1LmDc3DXznGtpB6a5PrdkH8juxDQB
3uXOU8FdbMFg1Qz4xykAQm68mUjo7PPmr39iqa1+FYmrdNm6S8ItEpDBp7FFaYCZACLEzKZAiSQF
r8/70Q1sY0eCgIr+AaSj2rkm0bz62Xx0O+QP9W3yqDO0Uo3zo75Ni0QceOprKjqgNrC3xYPhfyqx
TG2L8zksClqwKhwhgvTsddSo2oaeegQlsj2Q7B+z07sxUHnJX2l86VMKMudnCBeT8lKynxUYZqA4
/PgKF7CmywDXmYQnwm2PSn5GHcG2hVwvXQAjjy9DhCoL/jo3HAzt+C+yDJHTp/UjDgz3yrWEQYJM
+qawHZRr+ivVE/iKI4JzSShzoi5WNIt+65ohKw+LIPZKlgDMatEL+kQyQrV63Urg/l0+lQ3CPWsR
ofgDSx+83MZx11MWEtYhCctDlA1gYrlMw571a3jAxXfZ5A18zvpICkQ6HUpoEO5Tz8FHyga1+Gar
xh/ykQmii1SW86H72pKEgxHltVTWYotFlYq11R3u21yq7RT3WfDqiqCqM1PPSrUkWcmNq3rnITmS
n4LREV5Pgu144sBOWKmSvliVdblU0/xXEaxfN3RWgpiAw++aGRitMen8/bpBOiqO5GezWHeB6eF3
v/FdIJK1hfmUju2hRnxwpfDgYFVkDL1BaxKsaCOjQnRaJbd8bPXJNfI9/7sjUOozOKUNkOluGtnQ
8WLufHP8eP7A2JFMZgnDGL5Z518EOqiWSRrPlLVR2cNkLEB1sxh4b5fbLnPF9jhFovTRI1OBFvfi
vYvgdnNlOTzSVgorkSWGrqCkoczPozfCKLpqf+eVEV8RYzlzU5MyL9PZAvzA/rpq1biuKGCzOe4e
jpmqFUR05V4dyDEk/QLbMeioIRduWiSh4mtQ1EyaKsyArCBZ9ptjNdZE9xGyEFic35wvTcZjktSD
BvTKIhHB2uLIaHnNlG2aR3kdTcqLcvnQDax1AZ2A2RSPBOg2eFCdqYXSpUdV3kwkMDuIMaxR5e6u
bYI9wv4H0Wb29ovEb2lOY2QnS10C0/gMpXzSWjlrBfSV4z2uOzfSBY6oDE+NVVAwrMGO/0hALNFS
wvcEt8wPWQiqrQFnpujJpkXuAHcqc2qlgF8sul4LyRyVJ9mc6ibr4blb2qFi+rg4lNBsxYaheANZ
xEirgutzgcrjralMiSMucPdbS8lYcroyK9ACmxquYycSOeEz+AH3d+S8THchnjlKk2Mw+R39GSUk
ipnD3hiuTrZ0dYcipFxedAPgmiHmxFsiPI3TModKTvjUcjzetiMh8bZ6OnBaxrisOIqDwqi1vdTz
62ZBerOJAls+v+I0jT9Yp9ewN9dFCbfOQSTj3zwmea4d4PCC/+GRawsjf5TPCqILAOg1X/e3wyir
6WcVcLAuoDZJ7jGGaO0J2bEVzvCyo5nVc/8pMqDKOZ2aFfSZyVL+wIZU+gZ+fyw7kJg1nReSbBna
RRDf4mk0JOM6SvoeOrxaiV7WFdWpomRqqng3VXKKXHoEE++Flh0n5IB3hc4qzli45rfyl6ZaqFZZ
ssm+9epB2ncuhXIbCtmmUElGS5x+cK+FrmVc5OxjylizFzBwmE7EjSnOTFMYkrGXC62QoHQYLroL
tnw2gRMGZXGmDyLSDha18JGJRzlOv+Sh3tg9m8OeqSk8gZbHAgKAJRBeS0rz8rp06RPF1iCpjRGo
s9Novgc+at38AJK6DVDs+7xqjDVn1CXpW0hX03exC4CueZQkf8kVhsOWpbdBGOr6m+yrkfuzfAo7
k5Pp+vQMs42XyqWJt/aYpwqoZhX2oBTnCalNJLwUT4Fd3ceVF/1nktH7FElbXrlEzlv7j8J+Xl3H
rP4q0qNnGDXjpYIm8ViGU9eKwTAckKK0XA372T2OeFBwXbuXLN+ce0xSUJ+hdYxNvPkV+H/wbIdS
qWPQdz8x0VOwsBNWywguXzbI4ZIvBOt4U6jqY5JkbMEYh3RE70kXwk8ap+Qr6WYYpjNwALqug+J4
+3vNzyE1pDjPBBiGGuF/LwCidxHu2JwQlUX9CeQRNScbe45f6JtFWt2fwZ+Nuc+i1cfvcrPT7W9c
YaRIT7EreSNn+KhMByFVZY81WvnIt1Z1QVzDjRW7cANhs5zqilHnAYhCi+gJf1vWTLNKLNp0KZUH
jNI4Na5VzAyHIVpLioPQPJebGJDOu3bm0Yr7PJ7Jl2EEtk8SE5853zNNxbe6U4l0DCmv54c5Zrvb
E2airdvap0xxLtHGN3PpoytUv45yMkbY/PnbzitBNqsz/gm5kud9/1JwLCDW7MoEY+5Hob7aTbxe
hgvWuFGVMdvmprhMng58Jfmzib6XC6EpXE4sd+jvdptLOy5NYXpEAF0S6V0wO6+CvhBeOn5Jdpdd
dI8luz1s1hRZznZoJB3defcNdQoY8CqTssnTsYqtNzHMHkNQG++3wivOhYL9tHPxxy4SZh92qx5/
DEoLICOM+M0g3mYVwpjs0mtsU1+TLJv1Y0qThEB4DhNRsdah+qIELzFviev5sOtaBx0lQIg7wb7B
axakIN6FpyzGxZi7BzxLLZXR5vAQeIF/VNd4p7+gr+G8uXtpfX78aSY4yKe5mfDpcy0XQJIWFSOe
iH5lYkxg8YN7JWe7IQThVXaW+1KOkVxrUn354enwH7VJ5GRX0X9c/gzw5qvbeLcrwu+l61N0NzUg
N3sxdqjQ6o4UAwwM0pfuIJnK8NFngwclO2XlnQjchF2PM+2pX0G3bM0dL9VOXdwmrP8XooPDvFOU
LrH9kUhpzeFZik5REL+E1ueeJ3sdZEcafzWnhaNMAWVuSJJb2DI/5tiEhQvsfZGyukVZmzgwZ2WK
+sVxGr6m2OJ0Aek6unb7Xyg3kSEjIIxiatLMGh9R5dhRowcEfEpl6y+hFLV6YCfle1yQ23iC2AKY
udfVfAEiOCVEVOe42bfPP4fJ/aTRiEvJLoAjgh0OpgxRgAGYjUpV1PZ7S/Ddsk5apzk6Wtk+QsS3
NH5SQZxOBd210zZ4aIHfdiBRE8xZvrpD0cBqIfJ3ZUS3KEj7/Fa2bsRrhAQ+zDygA5cYKIZ1Vvzm
gyRyX8DLDQ5mX5Z2wUqfKJGo0HwqEazneERzxAQwiYnPCEsgsn9v3EUiOZ848Q6P92ewYto/n9Wn
IGVJMPfcgjaXb36168A6VMvVmQ6xIenUfL60VNuzB1FJxP6ueweQzo95W1up+b1cuEeRDKN5P/PS
4EjzCLtuno1V1/nDzVQHqYEUhL7dMoOOL5b6AE5dETEX6Q/ZgFKgynnlIvLLikt/sYjNTrS4VIs0
rp61zn+T3MmQC8IhYQ7akmqYIH/Z24ufzW8hdD3TwYk6ssplNSB0+A3OQWCPsdBzn1koXQLbJZVU
M/ax2kBHcCLepmADju0THa2zywSPDbBPTI1R+CssolQF4c24dZGBWgibr2IswNR3bTUHltAO80Lr
a8Y1voP37thKCIpNYFzCRKiSRv79XqnQcpt9phqN7VHLNrO0oFif2kbBzX6UKzUkzQ08CSME8612
76clDk67ASy5lcfsI0dHF8qcL45U6oaGvBqwvexum3P4007vQYz6iteqGDSfnVymL4Zkdgwdi40M
lCiJAFazq2AnKKe+ZqLkn59VB/tsjJPudoLy/AgmAy0qIAuer7mCmy24Gps0cATlhGdJqu0qM5Bt
lB4F3UrN4kWc2vA0bRRQ8CssZnDst5f0uT9eICV9quDT6KBTFo+Hiv2UONeEUFvHlG1y0aQ3KGhP
Q8VgioRj765KQbucTFRt5Wnpbm1Ev8s4xGnIRLcito6W/neoY6FU3fniN+wMESzxC785G48CzP/L
53kshLgovwR7LX8RRX9G7zMyybHsHMwjVOd9hXMArq7Jvh5bb4xQP6vDLb6cxif3ncgQAVz6sJuY
NukfD/nlpgJL5uTRk8QRxtP1rWUaBENZMzeYgpm7pIeL7zbgKKvl1IyrZVGWWc+ou8gRjXBplBKe
XjyxfEJw7ol8PwopFvcajJiaj89O6UlSgtkzjciLdq3w8IzWmX3r/MMHYv8BRgPklR4iCLE3R/1S
mrRdnHmu/BtyraVklYZO/X+t5PeNWKfJaBrXsoGEqyu/ObJAHrgR6j5KdGY41mmxekUkWRcV4t68
nmPlNFs9yomiva3sSAvDkTiPjKogEYsNEPUgrSiT6j2Pr7t8ZHLB2RP9JmF4hJ/xHi+ymNct6tIq
/LhmWL+QaVfmogNdQHHu1vfDPTu0rcil2q5HNQ92sMvW2TCYGZr6chIJyzxh55U8wIdB3MWFNguM
gEAJZIT3TZAVQm4CJqIf51aiK1V6FmaLsV0theR5xQqd1qmLxkkGkRBRRGkvOJtaFFtNouhKcje/
tLsUuR2VQ+1xvVy1yXNAeNfFuYsemNBQgYTRNpECAQFWNmAhHAsN2MA92p22vJdG2jr3nMNLBUTK
2xkeFPd1NetHUGLMwDWSp968ICxZzHMRpGdnvXZ8ECg4DuJoR+DLBcNaLi1qnm31AAW5RvhF9MqE
dRS3ooFZP2xTDDm2xrmhzRFBhQmr8jrZ+kFw2YKmNrKjeGNj07PudJNiHFiGi/giS4hIHdtSAuSx
4w58UoJtxE4iv1bbxiwvTHCwTutgbxBnMo4YZnwlEH37aiBNKwH52BgmSO4XTkXOueTp2Al7tj8f
Qvuot8DqOWc6pd3jKjauh2rzbU3bJsLwcw1rISP2p9qIdGj83v5Z9GqVG+bQG1VOoiSSDPBMZ431
3TpgVPweTW3Ui+Hrcla2OCFnlxeJXKWVlAFeFUgYupsXr85mReqKiGMGkNCni8LF65/whKKA4fwA
25ftY76x1dOkWzio1itwpCexd1GoYtkf6nGh4D05YcpaYV8XVMz4dy+mO/Q1XcLSSux40ax9FsEc
XfVBoOmGmDtkEz37yG3If8GEAlcCPBEzEaV2tPP0pEq6zfyDfffGqdMAb3jUl5Vf/TI0exezKtiO
kIZRb8wP4Xw7Imn9bkeoY4VJRYurcHNRd52MqTd2WAi7oegdGqh9sSHoFbx/060QQ+LfQFiVoCrM
OzXOf2n76mqCruuBjjKGYp1dJ0n+ev/B3iohA8qz5UI1Yxn3O0hGEoA0p3TpAYMgCfcvQ5ykjbWa
v98iOo8Y1EZYHB6cNi1hTH0j4sQlZOfS1Kb22dQNiQw7K+Uy/Xh0pJXOrkBxiU7K+ICnwPtSfJTl
28hYPd4W4AiCuwnuZcyKpudgDK9rKzXEfGX7JFRXKMiCCTW6vjC3rhQAvgnkdIyo82Mu2HXXA7LS
Kw4/f/Zj/wx3nOi1dEEDqsXIfaWezcwe7cnneVMIqQY9FLis8HmZAIrK/TNjiiAl7ooyrObpMFT9
dZbGVAHhu5GAtj1kbzpY73KEKF8kYA/bq9mfdlHq/tFn63n1LTTVROTwhNSlFb+ItMoJdpVkUOQx
v5CK/5Pfz0jEkEMKUZopgzTHDpy9AcTwU8XKnVtoeFZ4jMEcxNgQU99QwsqQa+BEY4VfyizTb92C
rza50sYCBFQMkJa2zXlepQi/p2pNY4PkRG7hU8erRKS1VeynAhHXsD653cq/jyu6biSFFi/joPPB
KlwRvCFsxgtXGdUzsyn85uzS4vSvBrcTzDkLKiTM6pIrAb9xpQUmQbT7qpDB+e01tmVtcKE3+NsU
gw/8s9D7Ddh7N3vK3qwwj43JYF0d62OoZKX9SOpzEmxtLQm33eNRoYHFERB76fQDLkf/2kPWiCS6
Wvrl1ZDktHACsc6G+yW5JZeXP2nMEnnT+xFY/It0pMN8fa5n9nQvZmwVIVj5nYkSvLWOOv8Fny4r
Ssq0XrlFEEsXNpviEmtvdu9YPcRfHXJW094Vo0ka9KUvmFLsGb7KtOfiEsux2Hhbx5WBPY5Cqhe1
wSkr+WXrmYjOCruAgOLAkezPA/Z6umGJs0yGIYRrXJjjYbJrF1ZWmPYMTDuxZLo48nX0wo4fxmkp
FmzWsKjOgB0/qYFOl4tTP2BmnwEXUCUUTbMsFAED83P1mCWEVAsU3fpCalCSpH3ZiMxMUORszF3C
3CGSgtczTDVo3Rq+UnFlxOghXEerpwqglkk34HrZD6D1kEYbReTSLPJZKTdFH95cJSYNOKoTf0OJ
77BBweLz/JOCaGje7ZtxjP9lhFXQfmXqK891/4yTArlMtqOK88Zwucfe+fOxHkaUZ+An/jcikymQ
I7zXoP9VvyI04VlByhW159TvkjtlTEpJlCCXHmf5yl9xTmcM5VUbp16CCC087pXUWAxZDGSXqqq0
fRzmldB/rKoyzSNriHpmFFFTMVPRn0kpyeG9IcFt3VXWPtv3l0Tf8FXGkOiOgD0xkMqEWVACWkM3
lGBulpvJl+Qv1B3OAvPlS/vVqTy2N7MTp3Vb30qneXEOd9/7BiR1tYvvtmUIWHWZzKgMl6xe7+V7
+1fSnfjYwHSd4AjjIjBimK1aNWHLBDbS2G2AlRtiw1gyWEWrnB7ex1Sfwc7zK1Njq8bFqIOSYRPT
POkR2SJ4R7sYGUEBNjrPfIJnjSjLE5/oy1iHNmo8cTyqwZeCksAdv7Q3HrJc+Fo1TEmHFSwwkVGS
aF0u1L2KSX/n2C9BpzyZuWJsog2JZ7MMq6oqoi7tn5CGYV8tTb0Cau8dhVz5OXMJU7kBFlUgAprp
GQMPGsKQyRc/UuPWNXFCyWG9atBHWBw6O4BBsSoQwTdzgkVi2hHxiiRD65gPkF8UsHFGCXNdjQOB
FVSdtIaQxwu/7tZPV7NeVpUXBvpiJyItEZLHVHvTodH5DDMF/Yx7wxpAJTTF6Lq3Ncd3ePG60mkM
SOkCbIJ2IuTjOWSe8M5Bafl3ElRkLkQoRhWgMEuEutRSLxRkoFUtlxzaAqEwqlQIin0UZEoJU6qb
x1vfY0HVsID9Iwa4Lc7aO9zkJAfQucoTtV4if1RCRtV4WnCHJ+WhVJXmv62jpaPfD0ON+2V5p9Oy
UeMsvowytmY8QZ70a41TErJA7ZBa4Nf/BnqHgl6u6B8TfhsLsF/fbG1aIO1byi/mNtENJiv18Mnd
EKSXllykoB7IgRaIzIE3defNxHX9r/m3pP1ACT1px8ptoe1kbBghCWks2ZcraNZJXbWvPkwuu7Ke
/9G7gNZuKy7+THhjqIlQM+1KjHOzmmn83D+R/ibVYqnprGNDTV1dmsf4NA+mu3kUMIT59UKYDHJx
hP9Ea1MmHINcO1TQvkIaU4i/rHba5qYGf+P+icLrdtre5ABHQ5GJLta9aRz6YcgK9CARmCKh4FiG
vZnA6mTODju/JzF0HRgKAGUQS9ZLYWERSkRvDeP6y3W5kMpJry5JKEfsvBJqTN9+FymyGW//9K0U
itty6WcIktfZG+PA3bwOuW5nOqVpTZ3mmMzXHsU8UVFMHXzq9wsoVRl4jUS5M5zN5VFXvFd26QCV
tAiC95qwHD3GlZ3ss1Fr7zhGNYICp2cMsGZSbA0ezT+B8iCd3nJssfsCa38o9RTaf47ike4d9X0o
ILREoYm7DLVIfCOw5ebTmR6nX08bMUJG2yiNfI4srBGVwxKU5Uc//etccZIUqZrZi2XNW+Qm1y6U
9yMx+k+uPG28j+sfzww6Fv07inFKBeYH10iXgqnaLVPtn6SKQ0Fk1PCthhuzIQDEUDc6fkVq96fx
pwF743gL9NwZDgmwFSB9Md5YNJV6CUZ/OBKNSPlI+WMGWtDCuzMfBfFepURPdEvMYUTksvC8HNtw
XkTY92Xh745jsDA3PUHeukM8fykmGuqhll6pY5sZBM5V+cdUh6HrzidGi4B9fi/4eKCA9D2BMgBK
aiZVDtonNHV/rHl9bmj8nvLG9i2tUCsI4ZJa5c34gOT6z7FFRj/8bzhNyYXLpafyMwBwugY4g9ze
+MOaq8UqB6YnNakMgljd84XHZQzFd0LkJMezil6gveYgh1Rprv8Mn4J0yDfYrtSnUKLYrcS1vPzW
iHKIpqf1+a5gGc29JgrQ8jzAS3RSAuA9izFaH+z7fgI6IgdqwQkW1/Yj5sv9dGgaMPblgCUR6E3C
g5f5XLdtS9vE4d0sPDHXr5YSs7ElEQ1FteMSsdhahpgGhHzUyCuuqucABv6BqXWfxbWHlISKW8BC
4TvSbD0EZhzTSy1G4xmROkZ/vtC7klINKZyzmPdjvAzYOH+owLgYHAYseoZ1HxRmtGwOqNQyQJd/
kd7kXVM1CCYPsMTRXNwZIPMQaljm5iADXrvhhC/Wolg11oodHWmCcHuIn26pIcZw90Cvf/k+vtut
74SAhnJ5qq1GCQw3Z9Aaz7QGhZ+S3472yg5CAGhJg/Ru5Z0vX/SOx1SMgJcfhXTrMh9uzW4IQbeO
iw2JlDcKZKF+KlFTT6fYIdQUpEoibcz/iwGUhO9nbOq4/xj8b5OLbVKfIvJXT2yodh4/a01ofISH
W6OAmWl9pFHKD2GernggULImLr67LUgnvZJ1vWJmXhlnRAJ2bjn0GJiecspG0+4iS307FsRSyy04
7Plj0nJ8rUX7BmXXWSl+nelJ7jJY1bT70c1lagC7OsBwu+RpUdBN+UX3eQarwV98ie5reI3QNiS/
WLLR0DdiT7ncaflmsx4ZC9nU8EunJ0XZ1Av+m/iDIXxBrAOXD1olIhZN0+tbUR+QN4/cKX1PnesK
DYWTk+Q2CusRuDm8Nywawoele0t+hD9qduDJg99xWdvzUFw8jG26h2q7dgnQ+O4rgAVtBJHl04GP
mTmFUY88WuWDyFnV35vdvmyxgIH9EcUsaGejgV94uFcIk3sRqymuTN/rb5sh36B7yry2ZMBkQNlC
D+eW0USnmqMMpFtjk7++I146IPvHIQ2V95u6HfHy4mW+JmzCP4Nk1EXIcUny8iZtP81t27aIzK9W
Cm79KFsWicDDwf59qbD8ZmBnFjUgMW85hFSya9r1ppcDdIISIlHHFnGxJ/7DW53KBIGNc7tgM7sc
boDkFzMzbdQk2wJDUl4sBZ7fFBSM1WnlYc1f3uorRxKkOiFg15s2Px8zYQwiwCwOaS8W+53yT4wQ
CW4C+8+/BFV2VsDUcHOMYj3jAwsWqaKW0MsGV5Gzuc+yzlQHORMqzal4JjsG2mN4hSRQnY9te5HW
n4xtyC70dpCzumK4o+I5KL8fnk8q79csoI+13CNd2jqeH10gDNnBWmJwI1NrscSJ8YS6b557I439
hpKjujdfqEPrrhV2R28E6kMTEq3WT7GLzLrDLzpAM3apToab6Nb0CWlkyiskmZ3UBYxdJeHxE37v
ctMfFEu6CYuWpXaf//IWySakmGyHw+I1xeedsUTvm/M4ju7YpduzSrlv3Jcn8ORAAtwF57SpHjLE
9NfAzyGTlcpYDhoThAPaxjKZf9i0KKfLYI+3tFYD99Yx/I6Dx9l6LcWhRUM5JB52Q/sorcPtLr0O
qTJYBKRfV3/5C/RRcDKs7nmiNUGiXSN3RaO+7bAx34h40CtIZ7Vf86zV60OUHnAb3Vtd0aYjZCad
ttt55YHWBE/kVZ5meSsyBRCCrUgvlAzYVruyHfOqV3/IgEa+D6dziWpnEjCGwKsrqFh0Dqn6E7og
dw2SBICHaxBo2tC9qs50f5gb0JTNiYYK0Hpldi8YF3lkP9zF7vlaeHSYJW0ZF/9c9jCB+7PjL6tD
LyrbLKqZtIFWJgimVYBox280v1OKWgqoBHhAy2wnf6yiTYAFN4m5zL6Hfow/VmroeeLQhSol7nHx
1JS/zI7JjpQiEu1NsdXxUsrbXEQj9GUvZGpa4ENLtArXYFGlLdUXkbUoAucXpSoNYmia3G7Y/F4o
des9HpE5Nblv9rgWA36Y9M+4HBryeDO1j/yvKUECxVuXpkCtLW0sn/GANzd02GUo/MyDV8aA+8Ej
MqByNseaRSiPnieIToMcUYJW6I+GObqn+lqm4K6UJ7/T3Tamo1YMhStpqvZSBHvfmbVJWWB0hWmJ
guw1gGFTCMbwSfV9M4QUPZqOjbSaa1XiS5uLGEc2O0F3+W26x6sPCpVvqGwOKcmzBVJ+agVr0Lj+
sxolRj5o8T1VgsZeCHUgFZDu/493pF/QJTwVaflusNvTYg8267XWVl6rRDXfk8egLnCfiNlRjxg0
dLvuxn/4beSEnDGYf+f1PALsKbEhTr+paqdjybsm80MSujiNfM5kdIiNIkh51f6UPfFV/iPt0/ca
0Wim0w0yzKlX7DILMvQoHEC5Vqb/fBu1XzMog+yswu9BdPa70mZyhMy2DnA1j6pW1sV08KXGkcTB
QL4qOFbODg35L+B3tSEav7HYaE32Uu/peoJoCk5cDO9JqHNV8yKGPGSnbiK4/hBGZ9qXVXLPd+ia
+YcEUFT6nHgnvBPdwHh10GO2joEc/xwKw3hbqOBv4QZuiqvEY5HWUZ1N6T3y+xY+Nmgs1rBujHc2
0vSMpyJdmQS39nH9NzL48Gc1SUFBfE1K6qXA2/hN85aElb04jw4BD40296vG/Cu3oSVN6Ui77H5K
v55/04BVMegv0pis0HaHnJljaOx19XfY9Uarhqc8tiLQlHC84JABkLFrtKnelqLdzLRNp8DK8YZk
K2lci6xKICymadQgyaTqZGWIBV95v7hLjst8eTbvLdyLqRJ58IH1nFd2+FMiLBWRaGuCJ0UiPlt9
gJiXATvkinaZQKtBWi5hBdAyoC1cU7dG1Px+qGTziiTecER/y7N0c0rH0CtJWmGyQ99ZpQLzNugF
46fzjFk3pDSpUqmk4Y+05/JD55uk1YaBXPI3Uvo1/XQtOwFY46aH27sVszfjKeDpGDa+dC4ngD28
9tj6LgqYCvaJ7xpWQ3QRnv5mgxUCk2xf5AgmEDSFD4gm/lCS2rPIe21ZH0RPfzhmOJNFYL/j+dFW
v/IQgP6/FKF3Q6XSTOjVUurfXBdxphrn0gXjCUzQSdwxnjwSVsQtbwUhCWw4VSqjPZaG45IXcM+L
cTBJCUR7rcBRPcZL0WhO7ADNR6fXNPQI35PFfXCZcUOIqLNMji8jueVya9s+4OpTf55R/6V2+odb
v1j8jKi2tfTxwDPXfMRS0cXG2H2rmsRyidCVs5OAPr8J+bhx8YDN/X+Gj0rtttfdOmhlOajaaOfU
3JinVFfqVUQdpiqnINmYygxBW9XcRExpEud66HLhOAa+bzDx5D3xW7kVdOldeWdZp7CqCVhMyGeB
k1dLL/LBNjAL665HEAgJTkT+TOCrH4snQJcZUD2TsWnZMNI/8LYh8OcWkoyW0baCbQKbO9P0A2/+
eQgp1Zru9xeOmcWf+rGPLZXbmxf4XlTMp7m0OWLxPw1OVdNokg3FwKh3gAR9+Rjhqd9Z1A6csOlL
C/YUOAp0MswM1QuW+/M+H4fUlkrbcUPQeaERDkLwpHKtWoHFt+V9alqP2I5YS3vR4ysWJxIKHLR2
/eWV/mXzUgo6FiSipxfvUf7L/Wk7+CtxxBGuMRQuMYunpgfUqQz9qBdCpS+TomvdF4+L8WEDVRKl
dFLZg6WWk7gtHdAzdJGABHoBQVymH67j4udscuSDPsfMFnuLUfYjfmK3qejQ5ZMfiKEHT9NjL8ej
uPKxfuQ6N34tTzGSUl58ayXVNfLfOn7fCefeVgYjG8ViWZ45ZHh75OJHa4vI+HbvWrsHknbd+JJw
IxFWUDI4MF0UlsFVvtko9PadOOZVGjZ5pUaDV1Ls+W2Sopz4UscaNmVn1dA09IlfY6eR3eKGisnw
BAROFxBdOLKg6CPL3SyD86Dn5cJNf3zr+BTu8522R6Vgu1ZEBwTqwJm1NNyxKidThj7SXsXD3Cem
v65C+ZdFlkvgBnkR30L9i32SlhE30/qL/FJhrCz06tMDS7/T8qjpmJDgP4XVFmmQe80iXyReCEQr
b3hEq+9iTnAurepMUKfUBx1QlIyD16w3YTA1qZyrtemLPS1Vh1Y5s6WG9E8pjvJeJm3GIl0w5o9m
l/HhR9TceCJ8aA4atP3cdKOphu427Zlq/zZqICz1HNFJ2qxA26SHoH8wRCbY/fmaCjTcl+zTCtCb
lpQyWOT/GGfdUEv1DGl53eQZu/Is7ehCXpACcqE2PR1ohDwdaps/o4vdD4ssnqZxGzVBZxUoXgpg
PwAlf0BhTMaWWLNq0RzyC2CSFf2nMiyN0Sh9TBEznzyyzxlEb/7w7oqRz7u9IPEJC2OSqKpYruIr
QLALIDhw06jSYl/kucaabiYNnxRqZDNJ4qPhQQdGZbERfmCCm5dN9f94rirMLwNIQbYnrBhr3QUf
4u5hrnNyOlWnD772BjJcR4v7ErJ+l1TfV3c0z8mnahsewePKu9pLC7Sng+9jIgHqfKHnV7MAfSMr
/q3W+ICCkcHWhuYYVdDXh5JY1nseVZiGQYZ1VIOl71tzdjeH2s/w9gOukuEUFMEX+WNv0WDvEWvN
EYN6G9a+/DT6hT9UyxRbjpJzMdEc8yBfvgUd8cDa7+UE0CpIvwrDmkSJTWwPQR9keFahiV1T/nDM
1HlHv91ypOdSFm+EsZ2kvtkIJu9GMXtXzt/UyfjA+W+04tHMqDzdidns+vetEXnk8QoCFXVOSmDR
4Gda2Tvef6GSTttpKnBSpLPwKuyM+/HSatUUKY4R0j0WhVkaU5HBg7UbdMqM+Wzkbu+6oJYSxyIz
bTgubGNQF2zvQvzCn1nePbrZJ3H7jyflnl4MovpiQPYshTVH5iEQzuVZdet+NRWVBcmNFStkjXxx
cC+mthIVRCdG8TJY4cfCBu2qs5ctP0nG6cnzPzItUo21uFyxacSbwJkxo/nbfeTThpVW5vt/28BR
HIxaA3W6ZolqW3zSqa9cejE+mTGKyEidyg88c8lhGSG9Rxhpt9WQHIzzwm9+eiHC0Wv2IZWQL6OD
Sfa63QT3jhRrwWzYNuNjpw2YV/LHJvtrMiIxbus2Wjk05ifpyyK6Rpq7cru3CopOJpbkekq+fIS7
4M6rLtgjRZLK2jMcG6cDZtprsIaYMCvykvacIoYUnOlQAs3sQlJ8uXPlucrsxmnp6YEvJuqvveP7
OB7msDPrtwLdjqc/1HxkqFGSRW7+JNlgsrgsU5BCPhAnS4M3gMMxdPuZEGuiZysRAc4jwHs1IrYZ
RWOOSg9rBYLF7DPGK1HFMsG+016NlyFskD+a/CB8pbEdX/Sndh0EeNDHc1G2TY9DxDf6itT14tC7
mpboEUEmbLbNTrgBl1/SQWdPeJMJWKs9haCcy52KRXFhBRvL5nMeRnyWPWwicSzsnnUVyT5QtjD0
nuvwgELTpGLZS3u91OVyqtk4MQrfP8G0CNHg9H1JfYFaPXd4Em0fv021KQS737JnLrFpieRBBCB3
SIbYKh4vNvb/NriMeFe0NOECZuJ3V+QDPNKY8CJOBNQk+NMpB8rgUbE1lb7wcuccosD1hjlDrGSx
E9lj41Yn9wERsK+U1Dq/A3dKG+TmnUwMqV2W91Y1/vSUDd+dUFtFdkBKs2En42d+wrRIfJKm64re
zl/7h7x9EQfcK5C2r8paNN8po6aLGwJhuiSkKa/HK9jrkri98N7P02eLW+23rVXchJQHiLJ7LF18
oMMJN8L0WQI9DlO8ZBmUc1xr9a+AZfqz/D6H6S+awLXDyg/eraD9MZnl7cTA1xB8MIrmTyjm5pMz
u43RdUpATjqj4TjGlNCtPDaVeDjYIxPHUehoWWBmU5CWuZImNQ6wghD38Ky5X6Pc2YW9OIHLvnM2
AhVDQfOhZoNTaoVkRtmJmsi1vkWEGvU6suqhQcM66jars1ShSmzvUcKAD7OTpEMxWPy5YwT4j4Cg
iYF16mwFtNugqNnSBQs1vxP1o4pFeaLv7NiHW/u3uz7ujOaybw+dILSOyoicLlpzETpH64kgiyoW
uO17tcBNz0TbbxX+FU1dX54+WwnRxsh3+xQbpEYaANoVrW2TUslVwCaIWw4yfmcmbV2AuukFfgIl
THkdlh/Dl2gALl5LB1E3xSEiTujByXTQ6+/ZnBsSGvB9uPg35l+CdIj1yjWL5M6oG4woFZJEgR0e
6j3ac26z5yfxTEOMLEvwjoh+NJggpv6wut+80jO1FnEVD3eLzgbDKdNf5mQhv86HOGWTEeTtJZrm
zHPqqDFE/7aG5Yh66vp8u13cY6emql2W56HHwZaGLTfP08q1rE8jgG6PTEOxMDI1JkXq1KYqlAiL
2zf41pVJL5AgA/8AN0C2PR8FvYr6jMYupybXJ+JmZKwPnD+Uph+vqZk2oqF4hUfStUcw4Rdjtxi4
V9zxnursBN7Gw0J590yqggliQV2dbNTHtArkTQs4Ee4VhxguPiUX6XS4QvIbJmOggEdVRDfUo/dV
NOSP0gG8ICnc6QCGU+MmyjBL4tvbxwQXQ6K4zgmUzVbklKtVAPc+Ge4p5m2KwvTz/sLI4aBcQHR6
26NUet01jPNe3IscekWzdsIHmrRWd9E3x+4MA3/Cea7f9OP1+TUvepNXh4O+E/nKlOnQrrBzYH0f
qSNxso9ZdwAdk2GjgOUK05zhsCqrI3rFjb/CdKVuCbm50QQlikWD+PffTi+5qlzuycn9Mb9hGuHs
dhycBxu5wZCvyj9iMJ2bTnaVBWLRGYXSZhHx/8uoM/gWNbFaFyJcOuLgVOW8P4AEi9c2UMOFou7R
R2tNZRHuGDvGZZxjAS72h0FEYNv2LmS+pNaJJc1X67QKckuRsjM3OC7TLjD6PVqCDyU3ycApEekD
x3UhAGdeRRt55V9hnshF9BBvWVRgAu5PkfZ+HNXB3pHLYwYT0QQDZZydHX3GZNok2HQ6SdkD++4n
OWUAiCCwJlm4cBfKFlK7hckfpN1I3cck5kyQwWMFomd5uIPirhHjXfTqRH7SJiANokXEz0fCK3vp
3iw7p6b0fLPaos4m/WgqduBQrMkWjO7Mc9fQBN2sL37bOpNs6XMO1/OgydKXRmZrS7NoN4YmC5iY
V2WPWUbGCpNa3GLwOWLNqmUvk8ayxT1obJ+ovDM9zfdh0G5Z+3vB62lBm4Azo02liZBykpHalC+u
TY2/BcL/3lCFD3E7CwDycIS1Zoo5hOf8PqGgbtqFeqYTSj3eZIXowoW3HAmqhfAO2hLxfhyWfCOG
VekqQxbmvpQ0vqs1ZtXQKfijtZsmzOt7FC9K/8PnJS1b3kIigtstaihAzHaLwWKVv3QD07raHx96
jkqs5zS2NDPfCNgVibAhEdd6YwvGb5ZYtDu5xmDZCIQmpIJKiWL4RZqzjt/URMmS7FpcrA+pAKGP
07XR4NhaihgbRBGTzyaWGOkvfK4PVizlfq+CxjPf72f4vveUnTP3LU2qWQsrqCNuZkEH3wHIP9nC
cofO1WdKlcSInyx6NXU59TWO3Ds4ZxggssBWD2Weo1lOrc+uw3eLWx+Io5/onPPODKRcngMJAbvi
oc29kop5lAbGv03F3Hkfs5xyFuTh0z96e05QJYwYNnQjJHwk2Jsw1P3WHpacrbecwPUkJTpflGhF
iyxcG1mWxPmooM9uEsAtoN7Ag8oZEDBooCqq/K1h541V3RffZcVqYAUTCsjO4+MAPxWjrUYllfuu
HxZLsmqcOYGk+JDPl3fD+VU+NylyvkyzvnC8XC2MIjLT4hp9iJ/SbF6UXij3pykVvLdfDk6zusRg
JBkt7X46qNK45ESQmHihkxnVN9w5h5bx+eGknhYvnMnCIy8vvC/8UFpSyNiimFr2DzI2AH8sybf+
ZT6M6+ZUsj65VItyPBBm0LS2XAEejAWnL5cI7vpesEyRW2vYMJuPJFz61VEfd0F/bk7kwTFCTOpN
0OqGZ4kZ/puc7+r9ZPJfyAvmeEF3/PffzrEr2dvr4FrafvKGS0Ikim91od7rDyRDCm/yBzr2xzBP
OVojyjN8M55+V7YPmnXZCQXhRP6CelTEYUKiEpAgAnyD/I+2C1rwojYgdMDXCo26G0hWuoM3RhIq
gRkT1LCPipeoIFU/fHajFMCcrw1ISouq94qX0uktaYodsTgNcDRPfWrsy6SfCIyvX13xgHObYlrr
1Rkh9qMbkm1eobLFOZQpW5Ie+Mhu+UT4IYjEWPFbC/xwvRh6HljyjmncetausArkhYKNv9PEW8WC
aqGJEpDJae1q8NQz73pQh7sIE04oA63hE/nRqZmDQJ5uvxTJRSQRsi3VRPU1NZ2NtLpOdj7cbLJs
ozEuQx+cSeeRyXDq4Lh7rBeYwy6rtVA4hK8XY4/apV+CQZ69Ow/yfaIQmgOg1BDUjxMH0Qm0HJ5T
8Zhe/IC6+PlvRHen86xGKOI2+IWKDWinnP2EZhHPUnQM1LBdchqtv8eo0pGtHQg3PyyDFWNVOY88
GcAhr4D/Piin+umH6BEP2/bH6Xp/fF849NESks7Yl0w8h7OhEehnWT7nADnTZj51Uwfrr6BfAlxR
oT0QXp9NgD34NzALRt8RmDbOUcCp4B9JZN2HrNuslRG/JzVTb0XmH5Tw4+29xeDQq9FEOu4/+n0t
m8UFd67fuDgJCDvtUXZLgDaP6/eHO8EUiuuPqVgKcNDz9lPb4/ibwoigsJY1O6Eh0N5e0RMExayc
JNzItWmxhfRL8ja3xFgS+c+RLkfkIe+onPBp+VrzHp1M5jQwvfQl8ktHU4ZDcyaaZ2EIT2I9+G4o
zb2x/danpsg5sZSjEUzDeKCCpJ34TFEd1rqFyO3/JLiUTUnjHSl3RgcVdzwjYAUDS/0vJgFgnSJY
WTwYDMiSAH1cRfSk4qa3160hPjQTPkA4uU4tlzrJKYC3cJ5fSjJaU+QodS78Ig1AyXlYFvoeM9+W
PN1JR39T3hR7KW/KPu0BWO28JbJBquWyaoBVUN9HWt4O0f6v3qE8TFT7ecFoLdTyaCMbxKXFVaPg
eNfHzbnd6Ch2elPIaNHwEeqlPPh4aR6JmTkv6rjLsFErBNNmsCfoZY0KQyFvNTNEJGEvN/Xkb9l2
+1J4+nV+SnKxrsoBpTgJxnhv9UUzXKRKqqm4YSmkm60OuDS8+WOHu5pjbPXq+mWEyMqeba8TvHFk
0rKDX1+3e0ulWeTzVhLWg/qMXcgnnq7hY4sEDBDRto4DnkSmVNluWF6bKmHZ/KK5rsccFXCwF/MG
vj0rRAg6Fyu+z8idYMTZjZ/+J+piphTw3hp8mOyjmpqBNjoJ/gy6NCLdmRxKwr9yjhPKNr7BWC6o
GC+PhGNqFsQ+uhGZA87Tmtl2QVULTao58jZQ3d7CQFttYorRyICyLrJGgn+Wazca+yvhJE9ORYcs
gsWf7yd58+RII6pIwuKkA4Lz/y0N0ar0zBLb+Am6Lo1htlWSZt5v5qacqytAIxgrnMfKpdpeIRWo
GLH22xwBvaljD9nNJ584pMMeguirubAVOpKuNNv0MNAFcYpkf4y2n3mSkHTcD/SNGWg/Uks8fskm
sLC8xzoTEv38ljHN+KMrKjhu+spshRbP21QkGSjEMHWoTTE9OZNLQQh8qZb2bsEL85NRor1IhmEU
0Ipis8MsSlzPqHaSyNI+fnvL4Np6JAsJMZUW8eRNuNEA7ILbRKWURawK/QAgA9Ip905OD99GbhsZ
wL2P7KyYZyeQL8lCCJYrZp14JVs0lThpRYXGi9msT2tbAikej4V2RdZM3R0UUkXdnH4vJaxn3hS9
UFCLHz9WZALUgCp1VXFZAb6TOOK13A21Ka5gKyFGEgpFy2mz14qt1Nm+cOjFu26aRF0YnI3/hOCe
MLzatCjgfa4B24WqMppHml2rcXvH9vceSceZT7ATIbdGQyJeTglDISst7nwjxDhyq/3vqchibHEw
Od3lwF3D8t9uAxB0cDScBjyoW0RoEdaf7iCw6zWkGp4/7M/FSoO1DdMQu8vemSaHc972VEtUDiZr
QL8DsWY925Dxv43wY+MCTusBd5u7KaDUuKGIOftHiAUjSLu6amylUPrm7u+ZaHjNNtkviN91dhIC
gMR2GEh5oeCbqpR0PWHqGtLquEnhIdiw40nvu/aHN4n0teyMwdMRV6e/MlRYqB0R7znJNZB9gjti
CnH17yE0WT3stFbxTZMhnYwy1CODGHOgcG/gfBtxrqHg3w++ktXILwxx+992c/jpnW0ed0jKjhGO
EvI/Sy61HOEF/zxw87Sbh5gj22A8YOtxp4+AHnr9MvT5ZROJ1PeymcY59IYzQnG+9vAtUYb1+ywW
zUzGPOCeWM2a1/MnFOXxKZo4IS9qpy8MROXzyhuOeOVopXQhWa+T8QaR9mRG59eaml61YjLDaovO
6mZ4dXS0+NCYqEKk0eOV/1u+BxXBsEcHhLCsQ5eiKvKQoLgp6eeElhcuUUpWr5qjo+x2vgCuiGjh
K/uyo7OkjXtX6l85v/EX2r+5Hr/92ytP3OPrl27nhzaJmD1BeKURJeFsw2vzJXxDz1cn6z2nE4Ur
Qyh4Z3D3qVHLBH4liMKpCHX0r9oljj2Qb/bRr5ywkAJ/PKr8AKKSIkGlQ5h0rsCrKc6WR25Zd7KJ
yI1y6BWRi2V/jZ9imVBcrAFaECLIhWNQUwW1LqsK3iw85889hx9H3+hOl/fge44Lj50FX7nddNyY
bt+puBimZ959w0amRW9lEZVOEx+IhvuVkcIcqzGvP8uSA9DxI7sdxKrMM9gVmF+2NAysyXvo+pvt
TZhnDGnePOsR4Pu48ltjABXbLd8cvSAi8A0ZTHAUpEcoae1S5IyLyFnUHo1p2g2lLMvZ1MBgPTv/
jKlzAt68/VPcAFjrClo5wwspKVpZ4cvXYPR3b2SswKO8nE2+hNlDwmb8jgP7AqWidcStGD+IqFCT
PrSELCiBSiphieORyL8Z0CtpN5vN0ciZWdVTPlJ//6p0ndnqHj2CbwlsGkJ5dT1436MqY64tBEE1
s4sFq/4lR+RkO/zLprqbNS7zz2tOsCkRJPioRxioK8RLUw2x/P3CIclqHWJQDJb3DuUc9NMTRFig
2RUj0bl2p7V4Oqlx7j3elHt4gfuuLTlm7P3RR2pDkrLfVdF8tXKHdOlbcawn7+cQ9C76DwGIX3qH
x9rjb+4dCj4cA1YOi+Vdanxlp1xFe9nyX+lZ0sG+qtWGWIUGbfn271agBkkroFlgLi2qIm8Atu6v
FOHXaO79XJmYE3Fy/vUKCcqqdTmDQNxPaaHVauSZNGv5WJiXskJt2il59bkn7YEXAc7sHUYZmVKn
m26ztIQT3HuObGbCkjqmSsIIvXyfvfBaN9l5+bLKsoj6dOfwbODcy+bVxrEAV0G31MyFl3w+prIK
T/WiYZoSnboUP/29tnzKq15T1cLRjUBGR5XntHiHmIh3U/NWyJo+JmbriM4Z5Da5nqouG2voDA/U
/4XAeI62/7Z9GUvjRP+yScnYLZRdIWM2lcKdjHSYOBuqNRl6e7yMWW8AzZWJTLalFN3xoDY1Ae26
+7kkb6sRNqSXQ9/tww1XVq8eGQZFS0tuIOhEsaSmZ+QBFy/urPvh2gFOolPFEcFjBKn6SxEpQqUz
81txoBR5m/ch69NQ49U+kO7ZZpi368ht7xWdoXPhaJtcHSdXNBvc4KT3gtg/gcEL+FNbZbXp8LA5
4szpW+EWaxRZ0IEoMquiw/4sXuL+wMaRClldqflVYgrRaht943JluaKwkJPNx0ElcUzg//9Ex8Nx
1xCWvDmDqU+nLPh0B/X6+5RYkm5FbOFFDoFbiCJFdScGqwKWjpOGcEP7KE6i51RAZjJCbb9o6UHv
5AbwE7Nztqb96OFxg2hgVFGL2N2ReSYA53hF1B2hGM8HHRLteXtSX5UBCgNO3CosHfJZBCWZe5t+
MJUAVGvrbQ3P6gnrviWrOgl6toJBEcjh/zHyrmub8UPisJMNhw+/Yj7fYDMw23x5BDetLkfpNeBv
nwwDKUUZ9eCcZ44leUrTqVaJBBF935yQrcZV4LuSFPNkJ+Vhst1i5elxqbr/UBO93XY3maSxpDzo
lsuzLLPZd92s9NoR3dqTGWYz6su8leefRKWW7OKvWxUQEvpWPHGhrIBwKaGPQwmdA/zA2gsh5tkG
WB8v8bX4Dt6vsuFc7tJFrFqr7tMsCAZyVqWGDADcf3jFbrS/MFV3m+C/yWLpMuWw39a4+rMl85xW
aQvKES6l7cy+w7ualh5kJL8lk6Vgkv7LcVfYlkaaaXOnLW5SEtb3OBQlXz/EY6OH2dc64y2j+e48
JmHOugdcYaenR30okVM3DqcNBQmfFwUTRT+qX0nHrTXLXcfkvM3lUnZzRKIApzvltjUhVBk/tUoc
AkbMJCB7LPHPcaIZ9h8KoiJmiKM94RAMRRZYqGuHNuL660F6P+oqfNfzfl22x1o5JkwpueGLGCwI
UcCRVVBr98ZsHC5yAOlZ6W++UqdPnwXRqA69CwHtpG3obtUZHlx2TLZUgUcQ1XKOJ7ui51kx1vTO
MBB+TP0uXl/TcrT60G3n1FGFdHg8sl1qB02cqbuRtwTxhokvTOnROBpwi/7WvYRpvnLX5taRu/pp
4/b6hBzBdq7HkPZjNetjKIMTnZHYchHGXwEEaeDfrlrF3fkkSryabHh/pc5XP8v7zHeMLaNzlVfd
upf6NR7a5rJjzR2CDWEo3zjlQgLCewNumTXZpOoEjnwgV4m7owsfq+rKVWS04WTNk/3HjpZlaZZj
59Ndd0+y6mxHoCLaHczSlW8fBEAp/M0GixwJx8T/jJq63iCAJxLwiJ+2cjNC8GWTT06xvgxlDIW8
Uo13smZWneRlUAToHEwP3o1W5sZc+o8fsVqtvHZJ57F0KNK4A0bvN0Vf34kWOOqTlgr3tA4bBuUH
P27GMJDxRMSkkOGsBgbmlRMaIKzbRdtMDihc4aLBuTOuG6Nsi7XxB7/e2HXse0U+jkwHBXfAARYf
8vypVl3U4l/AbsA+TxiKKCIK1Gn76We46xyGwKYYda4C5QHCfHdNLFkG7/8BUo3ckwinLG5KGYm7
R1P8BBxc/Cw6KtvL1iYy+TaLra5FUSn7nPysVDe48uy8AwI2US8jrMoUGjmZoGIZPHdRj06nchEP
9Hcv8J7uh/i+fbTotvvk6EYjWb827Kn3I6JUv3TLi4suZDnnl1ZMNyOjK0093Xs9nd5AphUP66o1
t9cY+L730+o03eIUMPkVqomZGJ1gU7aAV52esiZ/1IxTUPYcMs67lP4PYeD7N7QakFNduJ7ykAdd
hamkCmVB9qAxyrQXdTBdxm+SmiHuceQ2br0NqjqT4QD4/V5SU2guXV8+OIro52ezWm24aJLJ3cpQ
9ovp6ezMjf5yY3WXlAR95d+sDSsmq5d1st0dcWr6v4BWWpZa+Z3YLwjUUizb1PCKThSN2SiGpBrt
qGb5k1zmVQHcn7M3/caD4FN1kq/LLGxTUTygrXzbUN+eo21p221QQFgiTcABnjCFbAnRQpvFoo/D
X1Kijq0EdTivj0I692bpdnHPLsi5OBwd0cTtZVbsxJsAQFXQqojTirG4sxMVloJnELAlyFpjDa6B
2RtmHuoJC50bnOQXgPSDHDeFQ/PXQ32Lx3othzR9Cl6NVgd3JgziIjCCZ+ruVRqF5Kbvlo1kSRfD
lfurPmK/b4JZ/xq3IwqudNg8dZ+XyUpJd0MjdK2EwJC393MCD7AcsaoTk6daAoAcSnlN/hPG86rA
2zGCAWqZv4Rom7FDYCUNXVR04wX0gu3v7g6JfRZHTLSkCo4fOer44SGVvK1gqskQsp4nQUlBEudA
SBM0iVK6nLHJpp8iGzPIDGmoVuqS/b/4p8EqUH39uEiRw73GGIdUMT6eONH2gEbll3VoZcHdxRZw
epaeJxz9EAQedT7hLIHUSJesmTxSG9RrpbwXdvsOvhbskogjKQxvmzRP31kaSIwB8IjN+DK4oZbY
ik+KURj17G+lFjfiTgJm4xkZ4KQ9oWMhF8bNPhx71wToYKkdHaC7uPqKj9HQwN9X0MU3SC8he4iF
LNcLnZ+BHlGDFTrCceHsFIjW4G0crUDao4sIMICzttt2MKQcC6DbD/23bpzyZUvBi+WxK67QvPAP
grGzqsv0wIJ1a+DzZP6cjpaA7Bx47gEH80uULO2fHR9vg5J5e6HoiOc98a91Ysw4DGfZzxUGb06k
u7SlXLwoMXf1Z+lIDQjTK6CsYHNDgf/I7ps4aI+Vazl6bNZULWxTstVI9lQZprMH8C2KDh9PxLgf
VNY+6+sX+uOMnbZ09egPwTdFob6vvcgrVWiV9e5pvjWFqvz5N0XDxgmWVJYdv6N1XqHGtjtZ+NAr
a5XPonofoky1QgyWGQWO7gkBDBS0KOzXjXjDyeFbzRefdAoc0jzYcYhkQ2ZiPhehJVJCtpzYfPlM
3j78wVTZ0lTKB7Cco6Mw6z8Z79wUSs4EOou78WUdLT0dpHF+pGjfv+nv0j/87EBh4eFMjPW73BbU
09KhO6s1NyMLlaeDacp17qhTh5IiwPb16foqs8rtBZMIN8kln+9yb03WN3SMNXwWs98nGbKkqEu7
erfn+Xsn4UKa/hALsGigSJrJ7zKFAROrAfsPzHzPZCYUBWSqsaRnfD3XiTmqRzoNAgdUmKA6tBhN
X64EyAIVa8IDB/wCOqW1BFHYBUKb5Ce4op11XBhHG6Xafd1q1hIvdLvc+2/snNR0S9ylsEWtqXWs
ZGldFE0cTNscWqJTp33B9LSly4OqGfACbBYL9211UoNSDRn79+/BNVEDTcs0XiJJ9+zNr/IRr7cB
922w5SEqLsVYdc2jnyHm5GX2Zgso4cB41wVOkdZQqQJAQ+K3WnrbBFaaR5tgQL+H0RJH9aXlL31R
r7V3dUTtE4jjV97YGvc0PQyG8Zjq4Bd9t3yZU71Ym8ujMoAJvzixJD42cm5iIiKVzc9QUqGVmC9D
Fu8VKxCbHnmKCbsKdWZvjXfmzy+kOO/BY7hm600BiLkdHXZNTGsC2DRABLq30GJCjcFooA5KdNJI
t5E/+nr4Y469W6AR2vKyr6ifEO1YdnMeXvB5EYIGVWfqvQ6PH9O0/ytdwCSWETrvFrVe0MgpR7Kr
bs+k67QWIXuIx2jL86L7PSJpcW8Zzi7jQKhyn4/vkNg9YlFqeVlhVa33vy119Bn9P4p+/XlJJl2J
Na2iTb/GklpK1hYfly/5VvZBHgOR2pNMalU0/KMxBuvf8JYIcQbfRYkriy8kE5mcLfzrkBo2oeKB
ISm9TP4+9IpWwaCtNgRnEs5uYP/U+1rSsxNK4OhKH2Qi7K6+DJO+99s+n319nQC1EetrYacoVBjT
QPCKlb231JycA6LAZmafvN6SRI4se5SZEVhq6A98x60QkxdBEYQ2ao32InB34h53taiI0tXHHd0L
XOt3KapWf1BiYdObqSyaIVcJs65qGDZNP8BxKrFC2RLegJa3+M26FXhAcHiSfLNAkAGq/17pf7H3
P+Jj3/isROCL8xIVpAJF2zeCfQgTDJJtkWYhMFzoC/xDQaFyQnLxFhBJXarLGR3t9pTRd3uBV7PX
prVSvNbaA1owwBYWi+CLT7V+I823xeN9o+ROud32Tn7SGSSXF/eSykWhBJY3ymeK9Pao2rsKs0an
xMJVCV4qscvkQQg6y8qkTVooHJ9nrsp4+D/6BsbYj17f6thQZyyBXGLkiO++pHu1qdtpfY1yUDav
pKxC8wTHMCYsciOGVcyr3LozePaOxdTR5Y/IeCa31sAPu47ZoqMmP4/hi4QKOMO4WDQeG2KnxR/y
64omjhTPHyHyRKtkSjOZUQdNTwI16X52xTMJoOduWO83QDYpG7ZbC/sLFcREzEjMKiBT0xumvlVB
FVchgMDhoJPsVIPZ86LOGXxWyap3MSfrL144weObXsHHwQfA60BJqbuaWJccPXOM7QdenKCDKHVZ
ooors3FKhSo7lmgo3BgH5d4EC76fHxqOOUa9V6te7Fxp4E50mDFVsXpYoHGW+drNXCcIcBFKYaQu
+Pg9vFj+VBKOvVuRTs0QU7jRYOt3J+5OscQK7AA5UQerQAdEK2BG+NH/AQh2RSWguW43t+vHCh2z
dTU3Pwp5R4tn+UDIFENjugUN01Yr6dBQv/vUeULXRzWnSAG25C+4c74QFKWUj+P+zB5mnd0NK1jS
D2JWjfP8q9vDkJ5S7F9OseQUFaCceRH7l2llDE/IGjxiOQXw3Ga4eUOGXkQLLsCPAeciO0q7IEYK
jHc7faw4VxCYOpxG79NhYlz8Ywn+ejGrdX11dMQm+cx87OLs7Riwv1BP8Ps8hN67zT1x4h7e7/zx
wATgU97ViR17usTJtIPS7IcVrqjCsH621ZYOAuH6foPwFKRscriHrosEo7IIXWQwOvMdjD3lhtLy
9yVzYdzijtd6mhJMhjDLh5taGqYdJTEws2Ui+iB9AuGZbjBq2whKLvhifLEYtKVzXxp6gD/xrbHJ
SvWDdApf2pjNZ4iuUwAXRCrSvMBrC6CwbZ25VHXmz0ZokavN2Wxc+05tf8lR4xnAfzdm9qTuliNe
01lUqKeWwT7riWcyK5w9G+HN+5H17esavSsvFYdInmUSPuRgfDCPQOIpEK0vNAjt4nDwwNF4ej8c
dhTaYiNNHy+LVkqtCSrsWrw2DBvJiAkWEsGiPYNjy/cRAR8DYVKsMRNSrBWyx5vSYvXmU1j6UGtU
hxphCODg1JzOvu9BbSEyGTFHvFaT68SzdN+ic4ZU9OJpaWtsaNJzlj+q8Qay9cNK70nPbcA8+y+Y
DGaNIoOtZBG2y/m1XtgE4G4s0G6ylkVi5W3cy3iOzqXZ+Ktjrep6OJa9qb1mOFkkVCK/50a6XHB5
0lDGMUsAWf9zyJDwbSQsZKYpdHcRaohlz2BY2t78+xNOHKNQBro1VW0Tbe9aSoqfVH1k5om0Aa8G
NQ9mxk/vT1XmVLCYd8RutNeADDUszCRUTIVlzRmnY6V0QCXeOB38lRlOVc31ap8jPvPeT14xIUvg
s0wkkjl3hm3KgVmSsjJITxlKK4hg0VxGgf/+HjQHlbQoT3vmU76P7tIJVqRn9X9TeVk+032V7dJo
c3TO1hEkPnmXB0rKA7ejiXQoGhcXuUDyiuxRak8dlETt7xmVkjITMTa24g4tAfUQgrsuyIDToECh
IFBiFkpIZ7lFH8L/+x1Ju+SKTVRBEuU4lZcHE4CR2coDH9D9F4SxdHuL1iR6ZSM8Z9fgcXBt4EJJ
qOiRnu3v/OQBvzL5iISSWa76wblLM099DSzESY1vFGQk4p/7wG6GTtCKOyb22FC83rMwwmMLFfO8
JRNdR3NcVBqgi6Uo5my49HqVjjAl990YgED+dYyKTy85i4v16n/A6ph/XufgQCheGPRCcDTV8g6c
zlkLTGUDChzKpEKKtXS0SZoQsYDit//2i5ssf/wBSDqfdf5XDnnPsvJ/d/Ey6QFbOY/DIqhJZxzl
ZQ0h1bSucdWEXOv5C3tBZV+0x8Q9Mlx4li6UUU7AnWy2R1wsgZJLS/HuGfOQ09R3TACVXfzmMx/V
NFPCvmiPWumdVzW5s1Mt/Pud09+2hyGeQFGKlDnP03Dk4+k52Qp3ncCDaj4H7a43rnreSvrk37mN
uREPZ1gL3zA+sYVbT1sIew7cSpW2fh5aPilA9jIAuvWRHIUgPMwGcONgmthDRiksMZHrB3VTs5Yf
u5PgnTC0hTEzEc4viElWLKMFyJcvDgfeQj8QnFxeaVfoFlq/v0K7j4h//uS/8/bEOaKl8auP0urB
z7Y1xZyrNL2L9knwqTGpilWrPPzGqqfs8s0WdIa2ceMHeGoT3Aodg8sCuJZimJXXrYzBY8RmE5lG
rizysj6+pJo105+XG7DZZUd63CHJoisKgZB0fpQBYdbvSecmYWK08VU9Uax4nECZbwC+Frfbrrju
ImY8PCd9nov5rsgFQ8IUa+3kX0yCCDqVNnFHKLYFh4/dCEoH5ccKq3VyUgwP+9BLLzgqDUZKoFeW
lCRI/MW+CJIhsM/Ed5oxLJufUvUXMaCR1EASMMepk/VGzH0+CQPd58rJaAyCAfpmlkyoi3h0RR1f
D4m5PvjAUDldKmlV/HZY/EPHbLNJqbSXgDCGh2mZMHiBvzC6KsSOSTZIQF3gyKtqGmEIxwOfTx1T
Sc9HXeHMvcFQjwBRMMDnv9RQyxTcDWrGF/sy6fmBzlxCUsyHrXUhFZGphkg0zFD0uvk6OzzYk2BU
/28enGCXLxyLE0WT05l8To888ZXrwT3qL/sHDaqhNuJdlSsB8moVSrb76fPaxyi0ScZgGw9nD4T1
YmsAxKtRyFf1UABEU0CUm8LUqTKFS3Zy1MUmYHZqsEblbOy38TrSGXi+UlrIrswhXCpYLbphhOj3
UDc5iPpoN/8vjz6Qa+iXlWIk01hvEIcNXmXF6834aQdj2BLchuMNgwWRyF8aps+bY36b3OULoIwX
mnN3tvjQE91xa9i8CM+tI1BzhqOYS/7AouU/YrPkxEHC0WhArH8dpDElhqJ0Sl2SkSWOHiPeNEbb
BW8LJDaKBgMdHvnNbDIYgwG2+zXcw8Oe1k1nAtXIptd5cEuuek21n8vLWcwcCy67JwipXi/hPb/L
rSMx7nV+iPIASW1F4iuNFft6IAk4xWKjMF5fG8Ah9FWy6UXFzi7kT89neZPgr1i4xPqsDQgU56OM
WGPVVYo2R1HlNVXriA6LeZ9hxeJtCSBFpRtDnqJHfautHxDSYCFMAw55HgHaOxFsnWvEJtJy9KFM
0CPfCwcmBhRkRxuMqg43jVHs3VnpcWggC9ujpVlto/ReoYwCVgwJedosMF0I8e0Li27+dWEMKPt5
kpPmW/6J7AVmsUGFMmeB2Xc5NRGIsYCvupHyXW3ZBJCBGHm19Q9Mf46fJ8ut6w8lIWbNm+PsRY3r
6W7SV74tZtOgohvIzEE5+hJWKZYLbMAk7LBn511uIXd6TvIGInbIcb0wSXxYxHj4H1tnF92oBQog
vGYZPGbTKMSKL5sjmESCdLnJ1p+xyE2fgJrMR2JO8LWA3/mwrQYBBE0VY8Rtp5uZ4DFM+uSUhTi3
tS7DwvbAUblpCskV37YkS634aUim/VhaH0Hr/T5ifOy7HukLCssqiKgzpXC5qbhMPNTd0YUB6Ts6
aoB5+pQizQIb7X5frhitgpH93k7SbZ2ZmxMbYIZIlWKPqTR52k2Q3bZYgORiQKTrtIWCluV6gmW0
Ns2r3NI2Rd7QefPkX3Yvx/Wf3yvAfqtcTpDeCt/Acl68QRzd1FWRvt4PiljMd8FepXMo5bIt4DdZ
E4AokKx/mvYFx2I1dPVFn+yPDjISX6XtJ1EJB+zFXqrGmvNWrG6iIQUW0EIedaVORGqWVLzHaJsr
mLNKIo+n1IfVoWWoUmCt40oTG9rjfCYgffK0lJf2ZUv9pFofVS727bKfnzOlPeOG016YIZ+pTepi
q/zDCE51E0QhtL770imcVZSLNKxpkXJukS9Tzch9chbyEwW1ogRSmgoqoHbNn/iXtdyniArFCNM2
2zBTI6UQ/sIT6cWVWB8ly/qGl8Z9rlLtUeI9NJ5F9ey77OvuzCmR83eoqzjt+UEbQBAv8am4OC3X
hdIlu7HXe+0n/jIIjLY+qQf+aIlrXVCcwb1EjAI5J0Hng9211uwXTwhR4+SX9av1/WUHap5HB+4X
O9q57cCxLD4lp0qiyzvuoGZ6wF6sauFVjHvHX6dtvvMJjEhK/+uaLFfFCTBUeBTg5ZHZKxPwJUHV
KxnTjJbZcg1sIKe/PFh1aMmfkxFXzBusqAf76r8b1WaJ9JT2OaLUAQdEVmN3PNyPa1xf632ikthT
03I/lti5TXTpnWipp1Ck/jmISLGFJQ3NHYXKvzRZ9jb6/0gyC7x132i4vWgi2Y3Cm2F+KTXp9I88
wIL81uvf5fTl5LKFCI/IsCrH7Q31cvc6nib/0un/G7muFKDbeS+BEPP0z2RyEB0QHwmG8wN09Oe3
zgNTRL+BjIL+vebz9a7/Wk/thEMWILsQxcBm/meYQHZ1aMu2Ksd4vwjLx2Xjp3OIg2ZkugiwI2OT
lIzXSU2/F21hQnxc3NUwOrzuHvS7nckJtbX4mv3EKC+yLpZb4rEZczzmaU1Ickp509QOMyy7qfhx
0e8ve1w3ZG5sgjW4KRomea2yGRhJ73vuDUOuMprf/xvXSAuVQZeXIBDUY8rgwTFMxc8VXQhJd8gW
tPJoPxbRrBkaXN7sB6i9TinPzHvBsHTQruBtZv0IOjisZE7fiFi9CAG1IJN2sxI5HJc5bTESBWuf
Hd3oHOati2JYCLndBbc8BxhlT83wHWuyUXgwRfHdrp2kG8VyvXed9BjFowDmXhX2FvpEvtkgkPlp
U/tAj5aqZ434Fi4XM6Ul86FtdAmvm2STQT5hTlGoVANW2X/W8k45n+oXCE7tGhA5ojReUL0gFJgw
d+OFcJf5Vog8pUFt/am3Be1yG+LDraR5KzhSIb7XOHkcDg3CftAIutDzhrSn/oDjSRfEX0oM/pHq
1Udw0yLl34mWiYewt5E2QPRZVrXWj9Cfy2AmPbqScFclPOP2Dmf6RKGfNKsh89B7E82/vcYEz3La
o5ii36RsNGZoNRTqS7MpwLra/oNG1hfmkExJXlqUbuwDvZB6yw9hxFc4G39j6a4etOYJUina/mOT
qgWwK5I1rcRbe28bpxLb2BfxgG1B7K7kcmDeFGSDi+iKSeyqGVWiuyc7eD+JeAUx54I0WA0GmeF0
+0IC1OTmv+ZD7LEWE3xdFVENI5h/bnUM8OngstrWeXCYxH3gni3pGpeaR/So81kqdfrfh4a43/I2
3Vmrxdjp3JxxPuCBdgr4nurJTkVFIWyII2A9w8jc4DipmLzTXlBWcvei2fxdQww8EbqwiizpfLw/
xrabeCUC94P6vmfsucJ8F/sDj8bm0KnlVqjScxJte7/bjCF4jGJ1dyK+/quwrfUuzJD3+S8GXGQE
iFcGZr3PWnZ0n18VH3MjjePvlyOJfAMR5bs66K26PKC0R0b1lsrlefR/fF6Ks3D4Bim8ThM8kOjF
yny/oZKeT7HPMO662husixaTL7dIRuwgundCGIzbcZBvBUjSXfr71hA4kRKL2VWIOIQBYIrQFuyS
8JdoL0QP/afKcRpxLoQB4Ftko5c/zZPcfdRIVRpMNCtjDkqRlkkUB0PGjzJUVVgHtZx0NZgos5pq
8nyIyp6diixqukoOTJ//d17cEisJkylgdvD1Ie3ACZMLI6Q6hfRkUhtTn41FUJK0gIvh3uxdML9r
IamyoMAvvkB60wdb3heFflo63GzJvgAndrGUr4eB1GaiulXX+Gjsyx/5vLrz2olGVlKd5BASSPdx
fHLgNu8O4OQARSm3y2rozFMxQBbszpm3kRtwoiGvT1l3cxLIJ5I6mggMRf8sqtSecB9NwobiEWo4
XdXyvjibW+CVbwrELD1wSLXs/0nWcV4MnMQ1KKoMqTCogb+vvHPQSyZ5oGfVaL5mDHv7Z8wIu5n+
tFz4Nq5mArfVHUXcX2rLXyiMa2Mw5A5kyPNSD8DdXPBIQjgHS/H1SI/bhfvSxeYmUrllpPC9siOl
6EmqO88BY44eRxAeTOBOnep+KvJHUapcP+uIi94cHKBpP/92sK/NpzGqBCZbnQfzs26mhA9fXWQU
MjJQS8R/f9+bejzcfdaclyQqxKJPIjeAIHphlBYt08WRDKkZ7zHR6ikpogGm7h2miN3IhwXAWw87
/nCeLWxiy2RjXp8DGO/b/B17Wt9NKxiQsxF/z7SM6r4UXTByeasgPo04DM3S6dn91KCN23hrWSAI
WNF+WAVKeCreCqnxwpIO1You90snrDySAo3zW+Tb7BgpN4Uii+2dMfK98Edb+350kbDENMwmfDEc
lhVrnj7UyvQuJAkT020sgpQXMDsKzvTsClLlxoVQskkdaRKpg9M4O7d8miTs9/cUuB5wl8p2Ad9U
P6Y6xdyzkGwJlbPSeNfeQfzMDiEkDnPm/edLnxk6sgxNCKPqnjT5+QaAIwgcIHBM+aWtSv4P8mnT
HOq3eO9OH9QmXBuH2JDPMZEefI1tt16zVEvTmD1doyk7p72jmuTZ9NBBVC8Qr9tdoUEbRSIXPsLd
BxgNsmqfBq+PiLOX/9sarnSSZWWPul3XPOF80MlY6RjKnjo1+1G/zk+RB1+wQdg4oav7Rbx3Lx/X
+uGo51x8FXkCzRBWmIK6Yxgmj+Zmt0M3Jie8cLSGJFLItbYYFmnr5ovskbriweQ3aOR3waipVmhQ
aH+E7soLONCBkTybl+mkwfWAfQD+ATUO4J0rc415LYueTUigibEImEJrggF2+A1ISpXOk6WDBFGC
k3Dbd7jzDxmpfpvRafxivzYakrjN7MuG7uADspkd6g7vHeDxWzFXX2e5vFjmoZ8NrdY2eBlY2CtX
+AyVU9Vpq75pFS3t2WPSeklqafPdwskcvHAueEbuE5DuiDQEmB81ehokHlODrXS9zaPlbsOs0wwo
zVV4IKzwA5e4p7wJl4c+mEJvF5vSbfKnmwfDGpRxhpbJsJAkWk1yZABLmJ/xpKijEeNo+5NbsjAG
uDEaT23WvYbx8huPktcfmPxpqpw3LXbYZkUcdCygihlv5JrswK+tmKtD4jMbFRhsc5LNAsOoPo0q
G+73omgtWF8lCrhKQD6lWiMHso7nS99ipnzsH+vDmCbswOr2vhQj9LgDHpNV9qNX3YUIbZkFf+WK
LLRJt02RxLQam5dockCNrPsfHPLWChbEYajOBQ3HkKKqd163mbPMKnPXOsYeTBnaoq0U5JkYSPbK
y9JNUIl5lXQ+gJaq/FF8Y18qA/6q5OFRvtidDToSmHoUhQdDTQGNTQwERblvzsPyWmV4lWPfyHrF
uTR4UIjAHuO7RRAoRUCYBP7L1yVUuBpRpvniMCsSB6Fx2Tp07lD/6TAWV7/Q63PxoEnZ0VOwh6fn
iQnzS8EgU10tdLTJv2+9ts7laToKjy9rZD8bwRsPcLfyz+NCQOfvmO9NpZwsBFLXnWWXHiDgSLDb
L34MqTIB+X1B//Wle32TxFk9nTwSV6NbJd3eQOxuPvTI7OKIbZHI3+xfv2i1d/IdPBc3/A/04Dh5
TTJjxWf/EH9MJf5gWwV9cIXzkvC1YIw+5vvbDxQbmkhVX2Uql5PVMYHaO5HvuzgIhC6qYUM3DtRB
uE+kIR+337Y68QyE2KbfnjJjpbEhNwH2M6rFib/K4nyJ3OE4QQGYdY1DN3KVlR47jSP8d4xBTfAn
mgvF5DY4W3prLXpFSvK7rJYfrYifMV3lc7BjufIF65kz/p4TUbNGHbhMvsyt4UQs025E5AqbXI2+
jACkYkQ4bP+7NAtn6w9U8If4OCbXqi0GrcjKbKa8e9Psl5uKOasfR9qqiWkMbTtucOFFbxzhvmxc
hMtXkr1xREqufEUu38MzoiUn8PXcDPymUvav5Wg3CvEEM+AbzYpbHrvPjer4H2O/XvsTw9hkbjnu
pV5P/4kJYU8Gj+RjzIefi8/TYqRGwfNCE1VnNm2dUF9RWZevBhr4u7vr11sMjLyiDJEUhJfYabat
Ic0Myi7r1emaOG+5NYktc+4acwSX7dmaExvEulzDAb/1WtEYyEByfsWZ8IstMyRQ+w2xZYx1+R83
KA1aqp31RKcbDJdM10npKO1hdmRFPYwhwfCoajnhR+74TXp+6LAx7wBex8c/nEhTyxLj5ryvw087
Mo3kRZouKnfvl8PMjW2mDarXaYuK/H6VL16gwP8e6ai6K5TWypFC4sl1XIIo2FPSg/e7CcrWL6db
oSza6EDCFs1KH1X+Dvg8ssf4wq9BzdD96qlrVPiprgoGN6intzFfVXRTMB6HWtkuJl2J3oa5IeEm
w0cNDQlL2UVuoiuFY7GlI+zGtB7WXO0t3KZqKckR5AIL97mOUED5onocCYkCfKM3wFUMY7wNgNJp
y+As1ipkn602bKKJDzNEyvjb1bjGrZvttr+xMnaFV1xUIuuJJdE9QrUaoNYiar9ubCtihZuISDRA
Mf8mtFDXqnOYkWuVztoyzj5BY6jnJHY02txHmFORV7B2PlpdhDizFD7Emli0q7QJt5aET8Lb+vqb
sJWBGChjp0AZVj3NKxQIZrBA1RNDlUSca37idNsDL0s2r4/yMDkP7RPmLxgfJh3SFlHGiDYusbD7
f1urNIpGEPh0F7GBvoZ738eh7djBU/oOztICv3EqV10F3nIIA+LIfcvxTWpKFaXpn8n/de/kMpKI
pO6wGwH6bmwkj96+FvruZrUQo0/wnGxYhi2JLUGUbcVPsMbXU4pmd+9IYqCtX3ulVBcxuKzsPYNV
MNrG0Mm9Bve8PjGD6YEIFWnfz1uvEW9HClGEsiz8HBl066fCNJuplW0NTCmuVZVL5tX39Q3oBX1I
I/uCrMSSzOCIEP1/Qt/ijKii+o+tSr17/6AIkprkNprj8fy4x3HXgo7yP+ns802MtUCFJxhMtTb6
4ugkd8Kg9aIOyTPNOyHvZa5N1Lh8Ge8gCQArYF7t2KLQT4IgI/sDnSU2ckGk5zES0vlTEKUmyXU7
zcnqz3WdAasRF/f2sRjpABPBVKvpCicmkF2R5N2QhlkXvBqbMdw6wpeoGDNgCaNkg1wiLm8pRrxO
t9/41bwd+5/DzkhPqdLimYsiETN8w9yWfOYJsv4w342NxLwBzyfL7ke69sr9dwjZrG+5LCOrSZPU
PN55D5yhuAkhlERZLh20cbPPv0iBWNVmMEk+B3AAjAE4so2I/uW7KhZJe2FDSjkww+8QM6KvxRlH
B1CjN+X6Bq/keO3iJRFD8sKl2vE+sHyvjAMXhejvXR8RicGB3qN8ou/wQQryVQRGgM+znPVPEFC3
9UNbpfi5aazzhnlWXojE7qbyZDv1rfUCaPzLrbpxeT6ODqYLOe7V4FE08nBdgOKS3TZbyEQeU/Br
NzqtCLA7xqXK7QdMyt1+uRQyZWlrhePZfj8zRPDm3fC9tYw2vOMX2q5gFVUTciOT9KYyF6Hp0id3
36nydECK1slgHEQs9rxj5fMC/Zq8VHHEt4PAkCOx0iH1wY6I8wr5j7fwfepZP7XSF5zfh/6m8TYF
V4xsqkwuFa+r4jMd3zthmwx7Id7oqVY27f3bfVZvbvd1JD+XlH/kRxvqpkHJ7T9w4YD6mJpQza/1
XHPikA5AuJSy2t+aEUF67bHw/MljiL/PCqU/6ghYnA6RUNaI8gumtbJ/Bo5IGheYBy/QyEnA6I4w
piRyYaYzi87Yu79vchMbgIqG0KTZSX4JAL+oTAGnwfK7Qd/+fGkBwRxPOLFIdHe/NvSU6sOmhxnf
tVdVdPBzwX+SG5v2FICwXvIWauubvJcXxa9CcqA1UZBZDveGq5Z/ru86DZSZujqWtfN5V0BJEUl+
ua17sMGPpf2Gbjz3t/fmlsGLfeubyE7AzDQQ3E4xXlGUEXHlaRncpQYSbRTIbCQ4dMbbv27hMbzZ
qA8DMOSi6HaZH9HHsM0n8oaONrE4FRgE+JnAGkV1pVpmPSm+P0RBfzPwEheBK70L89OoGWmFSJuA
rQv3WegfdWUDJV7rWOYxhPdtKsukMJZ1A+fO7cQ5d7zUE7FkrLUVk5KA9N0qNPwaj2QvTyCNwr3Q
uxDNhvTMJNCTQsd8jZ/Yzt0SvP3lOuxueOZqiAtqDq/UZB7YXzclWOSLKDDJ1J3HG01uIOHy1eHP
WCC9heuWh5kn8D88uxFPqfdViD7jlSNqC29PyQ1fnV7J0mFG4Bgh2osN2ea5blOQE7eDfTZvITXu
ecmcXol3q+4h+aOOYDEkfyto5sT+zsN88GHistOQDxVdJJaljl2IsjxVA5GNY+16LmD6NX8ML2tf
eAWnR3tGWoA7mqPqSTEEU4TSheqHWnLFMneuIcIlm8twULWrFgPzecnyh3TkUxcnB2kKXM9cO250
r+WZjdcLitvPEriRWmLA+BwmhqzLv0u+a+z/ZRkaG18hwGbC+UeM3Wb5faZVPIG5IKJwW2j33gCV
32i7f4HzHoB4WYWsBgIbPQvMD8+5TOGwtX3BzxoVKsjNohhGYi5hMiOFMQjB/Gyalmiayr5CufJX
FxJ7r8eGenb9zxjGhSZkYMmuK8ztKiXR5FcElvhDnvAZZJstYc0df1oVTpY51nfYAB152X16RW43
MqYYZwVQ6cz8nhTLOPlhTjk7ppKCxKndqx1KB0mm2HOVqqAktdiKhwn6dhqGWboDk+/H56g8yYef
P9752D+d1phT8sfTNqlfTrvdfrw6lLQA7VFF5Yx6mS+nIM/x2DHf4rUwoj4S9yPyhdHOb54AVl4G
laYWuPLkP3wIjAZsbsutvKgFtJ+LeBXJUwkzCkn7cAaJSPV+mIdLuOs/cphaEnk4Kprk2y33dYde
ftaTLETWa73ENg0QyeAZrN14ap60GetJLU3uiFb6v4meVPolPNaxXC0PJsf5hF/zvsoEBURLmRDw
FPPNsDOTbMTo7GWlBVUdcGSnrufmXL0oVRE6BqeMDTQBQaZGTAPXGyjiR0OnGZo4mPuNjt+ivVD5
atC4cXGcfAOnPm0VTuk3EoVNBc1/ISwtnJsLuaJoA0o2xagjdqZ3fbCIxL3yA1q8t4IdDsldZ6+J
nWkZ4wvzXllT9weMNQUN8j9ezosX2QeTRj1YlUeS7F44T7xnvr4N63C9l07PFkITUmvb1IdFEx7k
TkzxaE6puOMNqcqdJsS3VIT4og4MaZMIofEwi+NvIsiZ3IP7O9NZzmrcVJBYNC9E2zF+V0eDqq0Y
sHbNKXR9VFETxRyDUMIyJaOijuKKYDCygST7syRtWwlyGBXSjZb7WLTz58HXqoO7kORUj5KcaGb1
toH0+DemX5Nsz1PWXNyZDNCtYeyNib+BPl8wvF8iEnhm4DZXJTWmFeuHD18eo+zpdHzwWB/pPsA9
E2LpND/rWIUtCRMH+oOW1nzXaYAfsTKbAJ03NKaNGtgDDkQmSawyWM/8mFEYes5l9ASrCHPlf/Nq
lQW+rH0NcumGlCs9/DrqCiw6OX1v9Vgwv2ORRX4xmIbWsP/JqvwIoJuSbQ80RDaN/msSBTN6IGV4
W3rbZgC3JSMe62TH2YlVznTH/Wb+V1G4yxDz+iVA6TCwUhTf7ZioLNFfZcYyK3TP2mgwAvOEaU5h
AUfAkslO8kpsCY9bEo0PwqLxRSvseGsAM2/SdEUOusTpKt/PfCMxLUtWeeE6jQUENo7QcutHyh6a
NMnLLtx2oToXJ41ENUWJEaOlm2LtcQgB/Rg78lWOI3TtE9xX8zfV6wUJ3ESFVIFXJ4pQXUjFAVlH
wlRTaDhSAmmxIT8aFgE6iXIdB+dM09U39lva03mA7SzfRFio53FKkwaVSA3vwCMfvmHTLru409bd
+J7akOjWPVPWKUmRvqupYdLnJwr8/TDCc8Ndpt4ZWGiU5FWeZpAKp3n6WWpUWh/JticoxM9DaGoV
0w00YXH7lqas4qK8B4TmzhkCh6KuDsEK9CdHpTGo9b1Z8Tr1056uPEDUSVvED5eb/NiELwx1AThD
DDadG0FZoVy0xC/P0DJxBrzZoIeJXX2bbfxIzER7c74UxO0NIX58Z1yWSpycj8F2ubYhdmvCQnTm
iG+RcmwZ1r7zBO19cPcNhr+7DcVr/ymhjfBekFfq0SMwwcPRb/6ElfuYj9hpgnXtc7XMZZK+Fol4
Z6criJ+YpRHWXFM2Y+aQ5RKgzX5PGe1SX7LNcfXb95ynoeap3kkMt2ETWMPg3+71Ws3a14PqbIWn
pxjOC2eZ94ULErqmNTT6xnkXoDV+JGqj4cVQSaL0XqXj+JtZjhvXhDIs1XvbX0nr3I0hxOEc3YIr
u6g+Hq9E1YVcELBJjRYDNzFuYwDtVzAZt3ztQasPrXhobpCnltH9PVSqobfY8tBFpPffh7FTKg8Y
MWUGWCvvrRrq5SE1VbkMkmFk9iKBMqS3nM/JlrVF1TLib62Ac0CUJS1hEQt4idEPMrC21Yv6rF47
ukdtECa6OIJnM8vGxNuhrqY8tCHDrJmbM0daTc7qXqsD1vrmRCk+Gx5dl7I9A8lPj71dVt530555
Z1Z+U580mRsppGKpvyAYeUiYGMuTIgnDrj8cDQZf7Xiq7YhRxAaJO2iqcxQmYqA1OIKrzQVsl+0i
HERpmJDWBy2IvfS8I7CxRDqbiiF/hJ8VlX6T34bWyz+9TxmVsenZy/pLY/ANjyafoA34vz2WKO3u
oiE8PCkFjNjwD7IAuauJc54uwLenyJNZgxQQG8oN19qEYrvZ4tuWefWE37GKtuwiVYO7HIDJ1RSq
5dEOzXDskBZes0qUtadUwojaViTRToV0pgQJdnWKR+oqUyC4fKo/PyQUQ7DtY0B3StcqfQ1bIHeK
lCY+p3ydTxiYK48DqoPLS8bmbqW9RrfU5DNSdWY9i4upNBXz1sfKc7R3G2BMQN9HRikDvGan3xe4
ZxrcYVHORiAhOUa/r/D9V9QGj27PcjBSvBGHFtou9+qBHGJLk+bSkkDyu+udNcb1Sn1ml12VeltC
ZR+kDtRoDDNPivtIaWRszngyVAv/ApVBG9go1NjmwpyyA39ZIwWHUaZFfTF4kSzeUtE7y+Q1rhIT
YTxqxht8veu8vY2DNSBo2l5N+MOEYukQ0CxNEElAhuwfsq9xzVNnaIlYzNcngWePyOWq/04u1Txz
YYS9OgbNZSSah6UGIXI2cvMdA/Qk8C4CCMF8TUiADAOlLaqgis7GnAr2qSY3XvA0w8xlxbjkjVRe
YYNtAOqmsd9v9y+PkMe4ED1a5W0QiWp4GQZcaA1OCbwvh+i8EX3ln0db5TuJpvlCHLBwDaG7+u9g
tU/SbZdsqBjnhGaMHc9E8tB0HWiUGhiw7ieAOxqk6C8JLiGRjIQs+l/L7Yzb43unEDuMQXnYadjl
BTl8FE5VuGXmw+dFdkYrGejhfWhrRCul1mDW+dDvhLThYXXnpd2y6z6y0taWMvk1IgOFnpBaNu0E
1sEQTiIhsZthiHdKqc12v2YkBbHPBupQu8S8I/24IP9xRvCTdE3KdfK8KK1Ssjp04jVj0IpLgjbV
wx61C1gdtn2fhDBE4oJCUgTz093ArDVJwvrCiVAaXZe/hpOHWT7h5qIl+InsxiHrzar+v74HDJe4
f4fdR+8/IyxIlYGnguobCaR7blviXyBWyjCYHl1Tswhr4bcbpNhatw4/vRIkwID0y/brR7/P3zrU
n3UPlGdff4lbeobhxOZ/V/wvT50f11+PCgfrrcqRSWQAgy70AgB7pjfxDEPdWF6+OLC9GODiQYn4
zXMYy1aBZRvGUeSTPQr2hPW4sofuHa8MLdofYlF2gZU5K4a9W+goF8izRW5UK7jaEnENo5VNvKEP
jLr6ub1ZBEpte22iLQ9HSjkyG7WS801skaUaqvjKdVHPLnMUPwBXF4yRlItcxAr3RgtqvuzFfobw
DQsZDPHJG/M7vP4o9S9fC5A3hpxoil4PHcmm3oKhbTNCtwTa42kYOMhnnSTBp0henAlO1G0/xz3e
jZXq9e0j7z/5g1NWFLlEeTzBPvMf9+Eeo2vM+cUoxywb8u9H06gYejtz+mO6CrLRoVSDjoP0cHnP
/6+XjnL8YljC7/MjTqkJzI/c4ptOMm8ITtTWPIz4Gc+9k1PSrvWzq3nR5Wq7A1UtabE6/HvUWefa
kp/rXIkv3rIjdA0fBrFBOlQxzsBD5Ul4tLp4ihvKF4W5wrj973svkBBIInAFl/LOkJYxj25k7F5A
cJIdr+G4MereOxdmq4HOADyy6z8/hmNQ9f/B7Gn50VQVA2id49sjQyPfjYCATDvy8F1vd7cUAz5x
LlpyNNCFpzi/BXY9GfzF5k4b4Fq6gmrjV0JQ1bTp4a8LIpi4tQGdDpvSsw98VLkhCTKzkrZmuims
IMDzCVsANILfMSvhQAw42CRyuWm3CtxsyocnaTyLixSd64opK8tmI3JKG15Is7BZu+kLyHwEbPIa
8ThYWWBTX7q8DioJTHGyMIKhBG3QA9cnv1pPXu9w8asopXEy6DHBaeS7d94cAWF8HGPPNno31zVi
fwZWVzjZof4advucEw9gKIE6uja7nbwKnJqlSL5jH4a7ysmUTMQ0gN5gYlPxOmMZxJsiulP6e8Lq
FNvM1ce8To7OUSdKGE23R+0U5hfestTVq+GsaqMXnZlb52O+7Ex84l2FH8pHHXkiV9Tu/KEDuP3T
zdCLg2nHN3aj58+A4Hlvaz4Etx9neCMeu67q946otRn+E75inyAuAztNRT/rzcQoO8ts0vYPl5TN
7M/YmRJeCeQSDGRAkT6Hui2Gx3luF1YtYjJBZamaIyl8RyzavXnfo/cy5cgG3j5J6ILMfrPzELD+
ePtL4bL/XV98ospTI3IM06eddqE9UBRgJygeceIQgv46fTh9anK1IZzzUBIoudXmlntJjz0qBQEk
oTVsHVN0RXKvNSZNf5Cl8lzfiPJUnJDQbBL/F5Elw6Ynehp9WFzl3DKM1RDn1SGDOgjTATr1nJqC
rIs1AIfnq7qTeLhkd0XJZuVgiSmnWTuDB3pbrImbkWJ0tjqB5eUttLa8ejRfdHktoE3wnzN94m7N
5sPx2KVrdClT0BKMuO1BFgUQMR8yfUqlwHrP81iydzdveKXa5Q1yl13cvtCi3/Bh/AKO6Fz8qS4i
w756OxKPKDsVX5rqYe5KPNtsYurefOJBK1L3lCJCSdGpAmbLtDZdto9nTNsAdpDFV1nVHLLNlxTy
BtPasw4Lw4hf7y9C/BK9vgnB9eZMiRl8JCcQsu8NLgSBbt1KgetQ/DGQO+AKt6Vr/uFvcRq2RKZE
+mPqGFJz8I5L0PKI5bp4LIxutnhjaNLFwBxNMG1pNcsFtk7esBwyWpZlk5uDfjSJGDXBUKfrLXcj
kp1W21rLpFUuSGFAzxPhQZ51fxMO0RChzEmK3EzXPQ+bkZb8XwN9pGkv0OgAOvyCJo3C4wNJl+EY
TEBrEwLNnYdStK3hVvP6wBTOPknw+ihs1ZPtcj2WflTAWJdHvMHkZJvCGMZbE5uDInj3dT1p6iN2
m9LsFm7O+ZpcU/q4qwIOvF6YUEgpaXtuudCBhTdjmRO0Ik88D7AWr9yYV6bkdahtSjujwsFhkhge
J4VWxMz+6czNlvvh2gEaHY4xcdgaOcIlv5ZsvMRV+Ai5qJ1ddD/3Vp1eLZKZ53fai4nDXiXO8w9P
PJHwlwAW6ip7XxMggoqJJQEZ68i/8FmCoQtDR79zfoVc4n/DOSoaDc28LFkND7SSeTZxOkMDiH+5
S6+/3yR3CgqsouvyYgv/evgrOgiYNu2BiXowksZ72VRj8LQxGeuHQM2FDvaFraX14sMUgZieUFX/
QsebGayIAnJFwO0wumTpGhI/wlPIOsomhc3NDxqX0Ixb6yswA1qdyyiMS4cgXCAAgj9KGOaEG7tp
nshWKc5gKEltEEiWVPSm8tSV+VNongwlj/7tRY+J+87VtXKHBdCUySlX4i8Vg2DhT8rhzSWPz/dq
6qaQKbcQ3gvcAFcgTjdVH3gYY3PUdoseV22xicgD5CqXaG+Utw9DkzVAlCGZZJBZoqXJGIIE2ytD
tfBpBVp74oqNQpt/lQM3EmbMtvyeIv8jiCX2t3WSmWIZjfN2eoe2znQDLhukhwz6CYsJBfagPc8A
LeSSPZQS2rpKVqNkEKi8tdfM0gTZw/C2zUt7Z0W0l9m2B+DV8FXq7YvGxvFrPv4S+AD8ky2qNbq9
MWOFhzPpkKo9XTKRs4OYASp8icpRLFOco2q5zQ2iQxG526yoJ2vy3HcZ0ey3RHMlTFyinKMixgfj
OhFMTBJzYCTfUVhKmLYVwTKl912vysQObgIMVja1zrMBM0S4VClxsNVvDesBmSkghAUPEhOgS5j+
NnVUNbcjr407s3CsBWbyyKEFOpk2Mdj5fDHIX/kodHi/MmswmLLPDaXWgnljaI7vRKxP2wiRgil+
9aOrprZrsEzPhxkfnZcnI2ho6H/NXQsNCdSelp7AsDTHs1ddHGho0S+Qk5fYljD4vjUpw46aqjFU
n12bxZ5ukV0hCqZ7u5VFGanb0vAmoJwGOt9cLX6dVyhFfzqLS5s5Oq+N5TYPY5UH/Did3jayDsBI
h0xHUFsowPFAVm7STj54zEB9VhngQdWqNl/GHzjaFU0PopBTnKadbT8vADgjA+rsg1zrwv/O8KHR
8XOPZc1rYJ1ZSLJll+pz4PJXTGnkluaw6o1epiaXGvyVTNOqf3J1lT7ZZOj+dZlddlxv23K4y9eo
xQSZgPLdfUnFgepMTxa2i95xs9JhG+vY1XiXx0fEz+4Uag//E/nE3oOThc/v8QXK5ReD1fBjqvVB
SCuqNPlwZGs7Djggi3Sn2LT5y0JZX7rgkHt+LnQWrOL8RMU7YkBZFlFcNcOUN7j3Z+GxeG/NLqfM
Pii/k/hW+1QFW8jH+p+ukQqF7X/nDwvgoPCDajazBZrkqBRc4wHjJpjkUalT5crTcE6YrB2sMCqf
/QI9O3sk5S+6zZUzfhoLphFbvoII1ufq/ycDoHXBZSSHJ8AFnsmccxqIbG88MMmHIJWFST3V3BXL
NQ7Jddcdd3rhx4YzylQyIrxb+CnMDWDvSY40cETdopzG897aHayNDacr1xJax9LhqUBYz24mbMTh
fYYrkKyu/dZRG0AiKw9+a+mG1cmpuTsbIDmpBBSA8LcX5357C6cvn+y+hYHTiNg7gBVP2+F5gPNh
Aqf+2n536C7CSsW8fFMjIWDP1MRVb78DHOKXxviyC5/c11HDMcDBK+LwWH7BWknpNqjn/S9c4dw5
APLfI2A0bNl8873A1vJD4fMKMUx8Rjm0KWX0pWv00DzG37j7krTn1MWP1WHZwPsjvH5fl0IpVy8k
zNtOxM9Ck6C6n6DJSqe+HFPe3SpejT2YwJKv3b4VaKj/HUiNpC1FuHuvHXKkmE3X8YfXEygKW0Hd
hoQ5AaQ1sM3vjmRKmwQsz+ddIV3wFf+sEP9u5BUo9bFc2/YXdWoXJIWNgShQlRqCbhseoNeCdAha
Fz4xHtRmQsdwyH/fvRo07LWUbftEoiMpzVf91chR++DP3SKLwB7OMBwh8hmIBPVJkisckTT4B/+x
eXcuXR5a8dcuwSZ6XPihQFed5M+iWH3dVW10bl1NDaP0VZLFsBZoIHbfsMKmgnKwyrNktt3K3NHZ
wAl8fUfcaqohC+4vanb31omJ+mDZgVeTke7sqVT38ZSkjlOZjCG3lHjHW/2XCXv3QZCck2GsLREC
9te9xXG7vL8XCHXnvAaYHXdjxYfogtblW0IHPlUKTYUi4q+0xvXqNXHLvOhZvMFTj5RwvVey5Ywr
wQkDN8//oHJb/WY4FAdSNTgXiRNYkVkTnjISTKvvP9mqBfofTS6y7kvmr3bDs9lstk1JIBhQUijx
Xr6Cbww+APgj1TGRbxdrzHS5Co4PKLmcNxXt5Fz+QrC+2KwPh1qxsTo71JGHGYScEKI63MWZuVwL
Gh3ZbBhI++z0ULXCQpkXWlmm/jiJg1CFvyw31HZAt5Hy5rXlb9pWPN/26nI7j8NDJnZgC9svtaL7
v25XlLXrVWjMCoDKbd1Z3JQ++SQqsIKpGCL6RaEeiFiWt8vDqD0/CPirDgkqgWd/y1PJ7l7fFRhZ
I7PqMpQzTNtckX7djKsPPRPjjYzs5MazhM+v9SU+NM8jCU1ATkYlIou9/CniI7OT7b/2ZCyn9ueY
Lf9fpZ3wh6Cp+RRyT5+KgHkHxfK+EkdhMuOqATBqoFzLFzszitN64IKuYz2Bss8Eoyv+59vfa6uz
6nRxZqsnnDl7SFhhjYCxufqUClcu5ugRZ4aOjmQk9ofe+haZ7i15++hFyKXn7YlofFP7aUWm0R+Y
GJ2R5x9Q/eJn3XPdSUcJRJjWIjITtTVVIKWFNND9dfswHhZcoc8Pzj0xOBBEuxUqdlvysaErquPr
dWEUvL4rre4Bx0Ysy9IgTE3rp/efcXHY/PgkVZYckrvBbA38PrCadeoSR0pXHypU/qRt6CPQcKvt
GLJDTG9JP8dYvtN2KEOna+NZ8NKJ7JtYnU9KWWC+HgiwqRncPnoKMWICIitiRb7zbJew+DU5tRol
t3vbJaogUTTFv1fntuj0EpxlNhxfK7Jo/ASK87Td3fJxRo3ih0hMKSk025ovnNzwTCCk4NmHJT2v
J6bWAASLor8aEZT3Cz0pMs5lD+5M1EqhH66WeOUsDonf9F2P4PfhAzlnRvbHR/tGfRg6S7SU8KNe
IzY4wXpz6AaAL1FhHOv5KkcZytsT5bl+/IoyWFA6FODjuz/HC3mzqVzUaeANNVRM3sonJ0FotDUx
8GmFlaQiEaWg2RJyuQe0bgJxguAXErW+tzqZbhftnkDUOa3re8gFE08y3EC3vczB2pFVlHBhjU8M
EjwXt6VNRMcgl2Qx7FYfdJR+IRNlC21xx9HWaxH/7y6U82uxdzMwciTMvjnk52QhbPRcths0a723
/iFL+KOygvjVH/F13BZpOEsQ98nKeOY5KB1JwpI+C75EhWHHy0wPCb5bAb+MEe/pVAaNYE1e8zUz
lGwtewhMlIijqI3kVZl+EqEEAf9py6hmm9zJIRvVdkPFx3kKqUQqwF2tIo28iJv/RsDmCS1uGCVR
n8EYZG0W0P6hlfHOlo3EJSbXyWafibh13nxINDfz2FbK3Ivm13K/R9zX59+7e6az1+NhWwWteUje
iAop5Q0eJYXCnyX9n9ZOdRDDmptBJAy5JPLiMwITPVlOug+oEDLk2oIhT9OXchfzOiVqzdhCaE8m
Dq+XtrQ/llxqPtAKM5FuaPdVrsMYCVn6M8S+0YEdwH67S2+oN0mo52NvTgU76Iz0UhBOcwZ8GR2T
SQYVkCLVa/gavZoIu9BUmsa1L6Eb3wR4o5MOBJ66Ogp8IJuvzC3VPrZD8cG9pKZB58lwIxVtf2ax
gAolvHjIbSdpxYT3hdY98DKVpU7uQ0BiNMeldObPLdAq4MY6XmzIHyhqU1FKMbm9c7yD2jfSjQxF
E5ugC2eyN/m5zuLoLgbnQIGEZ4ifuOwlfAG10161GzC0RlNkPGNsMTy8rHP+ZTeetSbfGnyZWAga
lbMM47dIujyFhS+dDaqiVj6errCHppA44vLrF39DZ0eDbx0mPxwwp56aePbBWmAJVm/SC9kC2LGp
d2ijEkzfh/I9cdi8BUs62wgTK2UncmiVZExpZDgwMK5F3IcvCJw0eE0o+mZiwtlFZ/DlXYNyCF3A
RSfFhhVoZiSMhLOEdMZkk6foWu12D4SUqHpvxf/IJQCfVGF0whM6giHfdCOh0QBvODEYLns4DX4N
js2i4azuwlPBKysmwajxjC1pwFU+cvWgGpGFiFl+qVjg9QnQaEUeUlD2R0LvYdsKoSl0Gwj5vzaj
nVVVPwS/mRPysFPxomibf4ladtuJrQBIP7pQCIKAfQIsdn45ug4CLzGz3xTRGdSrfklutRQgZsbk
a+zaDDpd5NDNNlg6jwl0Z++7su2JRccdoyfav1BW6SrZsWG51JI88Wl8XPODjeL0ruJ/DrxbpEc4
E2fYjFlWtERsjVcDfDfstJOBducl7RLHX4SQDPAsUuun5/qA86OonRXAyvJL6+ipaEgHzZsVMD7N
zVHglqWcTAGkr61BjfIvTzQG69GqAaaPPB6EcXqDSSzfyK0zNtQYe743avnaVbWewaqOwFIeTXLQ
4258Z15IpFWKvuqMaBEIrYD78vYYfcOBMDLujxTuz9NcKfpIXJPK+Y5KMhJlBzVzPhyuCnB+n45S
rHSt+v0QIa2pna7ypQBOCOvXmuDIuTY6yTnni3/cbdzAA7wVf+mtS9Nyf8w4yCxaFpFoKk4jsrW0
ZfVAOtdjawIeqnIa1JIKlvPt5GTYJEfgpmL2VggMvHY/wzKhUEPQcE5l7AIeZcAbyCjaKMS+Kd5b
JDrm4FdDWZebixBKx22aDKLm2WmBWfQlhmO5Tr8CE16Ih3rSwtjP4onRlB2Qt+e2shJJcGgBMPuK
RKHkjOj1kAA+VB2Z6ebTNpMbQZPicIT7GFsF945+QkM9oh4q3MzyuhzkVhmo6uxirpd7o8RjpRXZ
eBmBWRfCOcs7dL85XlwKUWEnHkC/4emN3gw0ap4Urdt8HKNeqG2YwajyXwVAa5VwjOJ6P1nmozW2
YaBYLuZPskhrfZ9+nDqpYR0m5aNDAIp9zdiPE/ggTSnOXDe0oxZPtBWux0LZ1DcEFstR4TJKX4gC
0tAIwWEzE8kJL/cPfMl+rTSUjcRq4LklTtsXIQrn1kxfSZ0qRsdo1gshBdnMJBJi25PtgrGQevgN
TKarPOFZVk4DjI/xLtjcIhW8HKkZPsIlT9S3bO5UNahjQewRX6cCKPBucH8uvmuf4JXQ6ydprC1E
HnwpWXbkBbdw18MISjaYGTI+uPtNyzlpTrCcybVsqqRmKJ6jGdhMFqdOhOoj8MCN13242yr+mPk+
tjvsKz1vVdV5UBagC08RY3w6+H7oyDPNVIPS2SrIwZ2qt9nGKHQpWrv67SLjNpQ8KiRHQwXz1hR1
XYKScPaSL1CqbfyaHS7WD5zHOdHKDVOQrRltAt3EDEFqyW2NgaEdgVcd+4OkQngL8IrZHe0s9I6/
sBLxVABcPM57BTOfwM6kb3ppEnaQZWC/eZGdlpq5ajCXvXwNBm/AmtQBRnYDqMFIOvL+WUGhxsvC
+FQSSOEnqi+9bawSEkYPPIQO89AvB/l9kNRJ5MFo+QJMrVC78Ti96xposs4hCcZwv4RB+pIPaDp5
MoaOiOPhe7WNT/hfmSlD+R1i7xjphrjnUBjqbOZIRkTrA8OEEqT9pQHHdQKBa1wlvhPxftyj9LHb
712kLqUtFFSPEC8DIdl+G1VrAXf0IHSlpRMn6/OUMIgSD7nRQ9Pxz2OZE3+EZPxxEY882vJhD4HE
6Z6SDSRjPV5s/R4el6rpCT4ZDQ9w7WvG5M9X3Sx4BClCVJfsQf0GqUNamTnn4j6M5oH0KudXfBIi
NYvsbK9AeR1+eEMPYmb/OLVlEX7aq2KWASL69tBx+HtHneLXV4PGTbyRIT6K96K4dK06KeQaAvGF
ueA1cwowFLWOSVXo0Pj3hruIhfSU3tItekM/cJYzh89nlNuNO51Acc7CV+6T3VVtc8lDX1q8svSf
wsG5xc6JmTRjF/V66sr49qNFIg94e49HOcwyz9s9Yqc1NGn7JvtOihaUTiqadR5ZMcXIZ8otZzuu
BtdP46UnbhFWfw87FgJLMXj2S0jlJxrtSL7sxxmg83n6BWzZtOqp7nyP+LZ/4KBcsimPnx9rWrS/
nOKpaq07bH1o0cOJJENl08fDJ3NFDE+C4u7VEQ1h0pB5ipY4kKxZuD/zqUAL1uLg0nYBHWt1Mo68
EMjLU49Flk/dULnXtO5f0TLaW3ATc5LCkd2zFYwrvdGH4vWRmavJWVByeJcHQ6oDO6jPxeDkDoRs
XiA0WWG71AkJ2WZJ7EusiO+k9KYfLEQHrd1BcAWGZt0+FqQ8V0tcrO5Wj0UMfANsXrEMapaDwL/t
WGHODgCVFJUoPK3fphgwSuDU52+EIpgfSfVJdPdl9eenPJineXFzD7Y3MiC69JUAmQjlx6EpFXgh
46eeDVOwvzPUE9FBPPQ4edbU7zh8E8ilu321za2jOiYQ3mVOxlw9kBDzjZH1H+92OkaMB6O9K3lZ
BGJLHnDiwhsUyC3Wwzl7oALcx2oaJBr4cfV1ZsuHTviSTaoDcXKXUhUjgw+8BhZBM7pTx5p4VYZJ
xqApkPJ9KE3hFx38DU+raC2/7Yl6vtLEC89XYbGHsjZVOXChVvPw5E+1lExFAh1sdmvQE/foJ27k
+/2L8viuhJj3TNhubHDXlyMhfDvJQdUqNe88ycVX4KWZVneYB+YPlQkGQX2eRpp/SeqdnBA4v3re
zW8EMZmGR7JAdGo02a6x4/4EY8iYFQpfD3rv4iAo7I41+TxzJEtFZUQp9Hhz5STI/MOnCfpvSV5v
BEVjZtrEJVN8wTZqlZzKvHI4IShq34xGvz7Cg82RgxN/NsNMeGwCH5d1uaBvCgy7S8F/z4fndujt
XeQc4f20R2uRDDew8awijjG+vybLPscDcviylkkKGcAwFECM36YqLJ7/2EH2M87vE2sr+pPv0JFg
ijrbecH/AI5Eh8+MQkCmsPw9e6b0/Ru90MJwdrB3fT2f3LHBDh0DDGVtDB0QS8RDggw1Qaq+Bdu+
73B6H8/O+6VFQy+aEhSqs4YeI7WmkeGiLIovlIIqmrnLdLp0br9le9elhs5qvKjSdKykNNNPbeVt
Q8/CW/Uyx6G52N6z//sTfgKF7heVZ2r49LLGjxMYDJkdm2QrujPGqojwTyOIKALbPLldiTu+uEjl
+OHwqf0tkv0p9Yon3VU80eINONKvM+ATWjQMJFKv+LrepC3kr0VRuLHwb2hQcPum90fgO+K+gw6l
D9ImVBk7EdQ0am8+2DZBXAHZk0LzEYW52eZnWwOarYMPBv6eMCMNT71mALEfbmJZLrLnOHbiN7hd
W6H1FGhHUW7bFDXi1KxD5Gcywq0n8tR85z5D8hpxcntNSML5IoZ91XZoufotvXnfQWYZft+KXiVJ
v4DohKOKQ23DvfEvkkiejEnoaevGPES2+55egC/ExfogJDc5JzcoWqT3V3cZYHYHNmPb8Szn5yWK
2WszY1gHC06NNofFCSEJSPktFr22UAmB108zGkcJGk3O+4RprYElEAJ8+01boy17v+a6xFlWDyRq
J74Vq4X+b4friVp4Y9daB6zttsOgf5jQ8lLyPnbJFEMg1wRPI+s0LeI4q/A8ORcu4SOvn2cpoOss
UTwEVvxxiQNrStja0PBo8FdBkZiYLAxJwg0AUBKjWUN8iXGbmDfV2tUwzFe4Oxw4vYwl8leh0UoA
Xa8c7eQT7NKlYZJf9Qh4cO4VdcDZ9a7QpDE3sk05LtrnzpjlazcVZkE5eYCg0xEEQ6FaRXKypZGs
0tnw10z0yF0g6IqEohGKNc6vSfjSX6DKEvt12SDi3UdgOU8JpmV2s3zSI+L6EiLSkjzVUaii3o4f
HEssI9ICMvyo7s6B7JvhdUctCo3QyFqN/iffrlV4t+4mHngyFhwMsY7/ekvRiMEdAJuMrUd9lsGX
OmrFLIiNg01izpEUOQYKSCwdL67SIOY9V8rMevBxGY/9+HzOw8Q1ZzF++HkED01CLGfBJxrHcRWf
eCK5Qc+sdLcHou9CbYkbL+IczRjby3AwrzJSSbmzsIAMGaIgQoHyCgQQxcD+8nJQJLYawCaZJzh7
nq+rJgSjpxMXevI1biBQV38QRfrpzEwx/A9EMg6OFae+j/RTSLSq4zRFJNcsi2UiyskGFreJm8at
FFX3GoJIWw9IDo4OaYBkQNfWI3prwcwl4riv/zOhVU2oXId919EGWZyXQkCHmZvNRV+i/XHvybIx
c4nvhaFo0KUUrYXrBZx4/HfzstSYqwE670+C68npd1HyUCAFQhRBCocN8ztBkGt4qSKwMggv25EX
vOtcOMXIOess/WBjMBOocdY7mZstarftA+KfYSAXrbEjjBD9C9400XESOU0psXjj702ZpA39/qnX
uYkELPmOcyd0IhFwIURtkUsBk2fwLeSeynF56cmj5AZuLcQAhRq4CS4d7ngwTUKXWTJmOpZJMURH
IjsQwxPOytgnuSWnYzYVf8E6pcJDGS4KsEEKfIokl5Gk388/zI2bGlYdL7PeJ24EXjRbMmvyt2cY
s8PLtLvEHVc7qBkbmVs24QYOa6GRqYoBM+OXEf9ga3+h/3QrCaPb2H757dpAL457KEa0bF16CCQG
2ef84Qg6RDOwR2GVoMZ5spn4LkryMFyVRqM15FJSNzVLmoafmOEYetMwNCqqZKViCbv1E3BLjw8a
5u6tcAoltCOfKAZXASP73Xa8H9aGdGKBY79cfVAOmr0az21thGxfgrlpbBWaacF0XuZfurF/TEBe
3xO2+oejpceV2NU3AMx5BtswqOng53Bv2truiBYc/sgFXwsoJNLCV2YwaT6oZxOKu7J9iNJRQDPk
TaVzWRtbEoaitHp7fNSkxYNPm9uZ7/dAtyzlJrikeuBswHf9zh9RTNqLIN0MN3nuhLyU4gJXkLYu
kSCuQVJgMYgT1w+WR5NSMJ5bKcCJMAvpo62sRe7OXrlq8IxuNxZtV5HxRdgjI+tWwrxRasihTBdc
ak9emxuA/gCIO8e5BoxVKL/63W+Pc3ju+oDRjTUi8+WwM57n4AbQE986/ZVQ8qaO3/WduS3GkiAC
D2ro4p3kRjcKNHe6iybOziJyXK+yIF3IwzOMSUTA0ftcvvHpcZ2wrSAwLpggfysG8pq/6IamumRk
Qu3GNtfOVhv3Re2tC72ssUojJlRryQ+VunErZq4O3yMSx+UZf8OIeay/g2c/QbvxSdIiMCIWLcQw
tvNCMICw/ktV3d/6YHDqf+r1uFIA70t/gt6kQr65t0tY3PnegLXEyqmDwi58mMbCTAzqMaIHq+mW
+ByWTz+1ODBwFhEAg9ZeSh1Z1VYQmahWJdDSwvhGuRwbI4wyvghEYsKlGV4da3/34DVqmjqbLQqw
U5VJtNbJH7csA0hym6i3tKNRRDG67KlBdAPpkY8/fkKSKLjl4dmfhv3r1J4vAGeR+znqDnILuCb8
uKc1VIxGv4GwBhLChfCaBxqbvOZwVcPFRfQP7jZOOiwNA8UBhA+r3pUoHymuu1jalZf8VSoqUnE7
13AmhcdwGjCjjxPXthAgHV/qXXMqd8qxgdfsqUA7A5mdKYOtcW4upy/wCeNK+oG2ZzmgsXLFoK28
EBpNCZcxV9tMGTA6t6CM3ceYawXCinkhZIN0Gqgps3lgPXoV6S2r+bKJQ+hElzBwG0t1IpxKKSXr
tSOjEV9vOBdf6jSCBT4JQ0mOUuH+OrS9cE81KxsG9SVWXaYAO6VeNsn7MgP/ajFg5BmltfyIrqZg
dkjVhkdpxqWW+lg0Gxbtl9m8VZjthF+d9cTdWbuj/C/JY5cZPthbQhzSfMB8yNx1WopNG2hNJ6LH
fmnyzDQ/ftmRWP0Y+B/ZxFC6c5s1wCPCIPCuiyC3wwwkeG9oue9BodBExPu+gZ/M0O8xbGLY8zoV
d2/FGPlnQ0Vz3TcrXRZLZoz3ab1UgiubMoJulCvwHGYZ0J/26Egh9IWp5bC4KLEvQSX+NzPzOjWt
pPy6JeWSDE7IWwajNU9NcRhfBlC0hXcsvRljrOHRNaRwhqEpgNqqT4fVlflaTER6SOd8Y9Fvrozs
ywgXkIr9dvq3VkRXSND0PpPKQtsgmz0KmAgL1ytYfto7YugxvWOoMjbszysZQg8h3hMTy6L90dNy
Pn2OfZV/704FMEobFb7OzkK9BVvzjyzbq4MVO+j7oZ6gAzvelzEe8iyLWxB8IDI+gARezaxLyCAP
k5RAKf6MnBYVp5xIAlVXg6RKgnOprITUKdauGvTPDo/EWgReAp43Rf4B82yFoRqANyBR8J5KMXeH
mnJudYyD3EYKnXLlNkh0U6N4TaGaxs9Z7bq1TB7O0ovDWpJRC6mtAqI03kcVh36hwyKnmvQDSqXO
Fs07hIc+P1PE+Xi1rRhxxI1pKvQ8X/xWy42spb+UNuw+1I3+0NpyFHAf5nphlbuPFZ0G1rVOKwxE
UeV4KKOJomvDIqr/XEI+lfXqm7o4jsvhtH3kN/GAmx9W744G/aF8fdscct0CooBJjJXWfIu/rlld
AGu5/t4G1ybzlbxYYX38uVxI4tdmYLlWC73YMunr4ekl9epxByWSOE2tAa5VV1lTTB5ertenYkI2
+k6azuf0/AmO0EKsHl3VDot4Vvy/JcYzAKAGDV3zQHzzK6oduDHb9TLWrFpYVSZhkjZqmoUAo11a
XT1KHrkJGKQdcea1emT+YKKShAW1uzJEtMPW28kzvwyE9lnDrMs5wxfbpSrEr13q9Q23dvSqFHZU
Ld4blfqEBaoT5/t4nz2paLbs6j0h1v9a9SdQTNEgBP4li1K7cGKX+IJmOs3g6h9R6+apYVo27qg8
a1jYo2EfZQ+g1a/B3eJk0o9OdZXIUaQhbNzHLu11A+8RXz+mfm9mf/drgzTtw2EgohUPLKjUTA5D
t49VxJIyvmAjdpgwJv0CYnPIWioksCU5za568OckzsoOqPynesAbxoaVzqbF89VjPEqYC+28X035
Y6YEh40wZWIp0iQYKTSzvoROBKX4NAUtzshd2wbSAF060olP4HQiCqwHPmaUMFY3xXXURoSpfMuJ
ZwJXAKbWwpw0fPYBQk+/sFA1ZUNluYwZTNQ2lV2wQSs9ek/SB7wteJpg0BLtjV/a+qBrIZqiQS9c
RsiXGjInyHKwfLAAwWSTD3u96md2qKj4YxkvNu//HSszkAUDGtH/4DPgi6co0HUiIKxXaAkb6PUL
x/iVUyKpgnW5FawUqFfs/mb7fjim5CYTiCXH2dm0B9UV9qGyYfSgXV5mrPS2Jy/9O19+hK0/DbsX
O+EmF5aMNkavQcedNE/aT8dRbbEkSJ3W0lZdbLNWbjLH/X85MgEz4h4BlY6+SZP70Ys3V6MpUGno
UMak08Uuv8uBPijIivrCVGdaZUJdTy7ZeIJ1g+E=
`pragma protect end_protected
