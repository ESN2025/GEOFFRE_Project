// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:25:49 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ox2uJ2infqeEfVIT0FBoix4zSnHL3BZkh9vVf9APBd5Ve3lsyatjo4FsdTmnCBGK
Q0Lxljd6EmODMKt2K6pp8msIXn9+C5qGyugMLmywhm8MFbyMhVMihRbgA4yPJOp0
ZAma4FlZmadxfjMv5ZiV6lXu8u492oy0fP90LEIPwnc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17984)
AhbkEwUzOLhBgFAYn7oqov64nTXSFomV78fQuYy908T66+GwB4BdNxNXi3fdqI5S
jccqnmyyP/ojyGK10eUdO5tbEYOrNEcGOJadNmmrpQu+f8HUTL9eC96rBlyhC/be
8/NEIaD8R4X6p1U3ofLNwBcuKmMueGS/3tLmBOtI6ucDCaDaneJ+GF5hNgfx2tuy
xtxUVyfdn317NLcsncMHn35QxnHEbUs+5Mu6MnxaXS3uDHA8f6mB86QoL4kfox3d
OEDWrYmGjMpRQYk6ut0grsXzis1unEXJAuGlrTX7iKZDAJPmBj2C6+0Ccr1Vt7uh
rfLGG2UqJsF0btRWUPHL2hU2rXyCJLbtRhSqLx7o5I3vsQYV0eRjmT1D+gsa/6hQ
6mS6PF6S3wZzZHIZlPcAfU8+ONk+W+AkHbjANO4NybSLOUUSUv0GFxxKjZaHHXQO
yoHbNHLQri1qVuQrYwaJpSBRDadWZtbSYacdLK+X+qppJfxJNTK82/Ta2eQZHbvf
f/P6oRrm8mc03+BdD2CjVY76uDvBR4SiyscIVVYtTvL/1OkVW7RDy5W+gmRo3RyS
9T+HGSy3W44gprKF08KbKXfuDxw0iDRUiW/MjhEf9mMRG9J2IyLBGaQ7QtTa4SyL
hbV44ENvrrnPIIe/M29e5wuLXWKUi5hR09sjJvDfa23ve/WQLIUbTYYfY+WSmkaY
Xznof/YoCI2sYzbN3tTnogOAJsxYwNqeCFp8+B8lm4tGhjo8hhDAdpEsq3po7I1D
Znthmh5P8rltguZOqhTUI6wJU18TnQSfaYMZO7ferfqHV7eTyJBaZetm1eMRLQa3
RzUx11V1ghp/tmj2ib3Vus8pdJtMpzEGWysKTrgE3xAEgFZah3+1dAcvWmkw6JGN
cpk+s6uBh6h+bYgvSq1xqheQhOdkMdc3fpS2U7zBRp/rV3Otkc5e0uIUrhyKuou3
A8JnXyrem61RTm3m/yEMrNiOgdxIanrS0NM2Z3tE0PW4uE14BtjmXtMu+7E+iXCJ
PJju7k79R3l0VPao4fdd1YQLIrS8DDzOM2R4VilTcPhK86ScdHS6Gy42/ZVQWbcZ
O+tpBmSiyPMA82fCI+RV60NOURpEVOZuFTbYJadqfCCanNx+Alni6Kr+/n7+1QNX
xdOjQdIQ+09bkUDPgaKiTGc6pCNJelLPVra15bAEida22pEO0EHAGka8SVoWfxfl
KlqSrpZ96E3j91JnPL7+YXlzjSoyAnQ6C5MAhL7csOvdmM4XLvcYc+rWL2ZTseO4
fPmcTA5EA8p5p/39ToV7/MA652ojCngluadWfO+j212jpvo0J6mTrA9S0bBEt6hY
b9BQ3S2YCTNw9SMwrIPlwT67na4wRWnTrpd3KeibWfa6yleiaATTLPLLTiwfEycg
22d2W4b8th538oF18AthdzwJvmlkk4UMo6C8+XEEOu4j9xoOK+Jj9ExmN2z6EYme
i5T/vCvepHxtjW7q5oItotEuld5NxadMlTSwvDVRyWQ0HqBt9+/+HfZ3mXzxUQ91
sRIUKWSektbi9ZG+ENeLFzD5EuK8HuYKHiGPBgAZAt7P2l5Rspi+xn6N87ULAgon
0LoP4YL6UaTilC/qlzbg93HrLtWRpefNUnECLXf11URS2GSzwx0XMw0nDpoTTE6K
ogM0/0/HH9lFKU/6DQ1oN7Tn7BIyqJXnLeWBG7CACBev4HM+O5H2xZ3CmIG2G//Z
oZhgDYHUTKFQQx7D2Atw4p/rfYr/A0qECJNhRVIfFnjAl8ZdTFP9Ey7yYdDSIpcm
5brV8pIhr1lBf+RFvcEwgMnv2Pe/KFkQTNLWn5bmXZOBruAZ8c2gX9csynWqqOdB
6X7b1pp+GtsgNwVjhVhTZ9CBqf/ykMco7WwBM1w3eftWAia4x/WZVBDTSJz07jIa
nGObhDAARDxwj5BXuCt2TriCdZIlf/+xnaTMv1FeqPX93RilsSQcdl4qQVEJcgI3
EpWtX1/EXigGyV93E7alHxhe70fK/ie1vjFmkLI3yDb9MqcjVSRgDhJarNhJ1ecS
7x5Bk1JNWyyTH/FeEO2ARMP8DNx/HikIpPYsjEi6hYKtj+c7TRFvvPuRkEB7IcPa
v9JrH6acy/KuME/xWdlrNLQd1I8FUfpUzcKaa1QOkTJjHGk9FAoby6F1t4590C9A
YaVpSvBHRfbCrxS3dyCAw2G0tQ0rUFCP6HecBVBDzkWkCH6uN2BOGcCGX2Iy4keN
DC0xC3Ayoe9RXs95WTymGTVLBHS5+ZtMEJ0smC2WeQyCeSWsDzs3xKYeCUn+NWI4
JTwfyjMrvnk2qUpAUT6bbJGHK3EI1f2kpn+OUbk/OmnOR0Lr8xkmKvxamT+qAt+G
zKpyINJgY3vIzlrG3iWKy7/hyrU6NaMYdYc1LWKoVC8APpjn3xAAAC7UoHUeVQKA
mO3UX9EUIOcOZtBcv/q+5A4N1uInsFpVIM9iOhalqWMsai8iiLnJggGSl2HVYyGt
XcPDzhhX3kIhWUgmrVo7r0dr/KoyZaZ+dFbB9iaPEcGNWYTqcLjXC8tYfM4gRiAt
wOOBZS4jLNHAEPjZKqlf46AjNTpeTNS2BY2LKoFig0XfzdrRlD2TcMU2lC1+aV8M
4l2XIjOaCg2tHXzoRKlhw/+QPorTxcCA7h7YfnZrykkd6j5a1grF2L21WZ0qkgpm
7vilEiaTVBHMwjKZ1HRW6vD/jQb/aXR/0zdfJbRy5tEnq9w8Q8WOK4uPthVqFhty
c/AfRWIyYsYHq+VyBm0tNBDc57t1n7ODVT8PJaEw5Uv3Sq4MkOLWyuc5k7zAbxA+
w/VaE3oASJOxWxINpIkCsYZTTShD+q0QSWtqR3sQubkWbsuLsNu8PEqI/xrHEje+
h6BDXAL4o85tHEezblctDKLQersqfO8W6DCdFRpI8967t9VP8aXBkqLSBV+mZ1JT
U5xUuQNBlLY8jpAFykF9wE33E+dUjwc05AygQPU2IPX1NTLNVqKkZJ0SdEPpPymI
Zo2qCN6DABvYY5c6gi4VQzmcgGmrcW3kgpoBNZhi11F0g+pTqShmivkf3+z+C7NS
fyqVd3zfqX/2Ob32CwEj9Jy0QqYg6rTyqeBcrzETLoL0mIVOOU7YUIeSA2EQ/vve
xGeOWeIxOkX69jGLPK8dgMhpIVBS/pPXmbdpogo4lA2dnrAfZmWUrfxfTujx3AHi
NDf7NC8WiMn4m+w7NoeEnuxARIKLBC8i/q0/w3fbdcUoirltwUzjJsOV1Nw91/Bv
W1TXHNCvEPiDdtR03oUN+Ys+CdgjZF7YaTgaFyla9zrivTuJwAHqZ0BZV0LVze1s
mgAXcqsYOueGLi/15IOmvWfnUSs7I95/BbsS0bYhAOx0VoQZKJcAkwLuZkFUCC+Z
mWLUmVIdZovEaZiZbc4OJiDtJ10DFIP4d9iy2X9s5GftsAJfggUN3rICaUauvOfU
saIvjakFaoPPuMjjTt8Qet1fZQMR2ONw/tPMy5lNBZJDt3cVFIOWEirU+0JMObuZ
IXWMIK8PLPYI1ynyRmM5UXMGW4FI6sAqdkZgzeNicMpmIaOGDfLHmsuTqSRVfEie
tbbVTjqykaUhWc4IFGtSjGtMADl9Znvx7Bk3JnnBykRrAVoZVg5g3dOScVfb7K9J
wFBanO7QAZaAUXQtLfp1/jadXUGpTQSx05iR/wxdkDpFuj1uInreJ7S2WE+zbYfD
a/u+wU+oO/UzWRYzO3llNLQr2O4DWrcTy+xW67X9Tn9hZAjCTW2q4EQZn3hLMEZE
KR5gQQg/RIzMrg/T+5zpzNh6OXnRhFnhqH7yOEqHgxS/7EDztZzioU4a3zCnQCPu
NZ4So53PWEGDnz2mrSmUGtFJy2gWQRlICUPW2NBWFnhPq6Tg12mcBkTICZBK3lcX
Am/0frgojPNnP995B0naVrqYUb7jLAhYo0LO1/K7ZdBAx3PgW0OkanUXhYxMWbRQ
saDMpAeXcB+EoFRZODIagK0hwL5O9dkFtGUNiz+6hdfq7RPhraULfnJ0e2Tq1mx4
AZfelAHIX6gmV8MOLJzXAMDIjQfFiUhzOSD0tX9R+dID58axllsGXSk7K7ohto06
TQ2PnO5RCNRO4duijn2E9fZLFrYp6/6ivZ5CjhAednaamWtq0+bgmAdw2ux3ofVn
qmIbWGDKd/ZLH2Vp3OxScYFGFdmDZm8kjnbut+lJrpEVX1Pq8BvGRaC+ukqGTr4R
2f8dehgRJAnsmXoUWJgx+AsEAfqjYaGmdu7pHT9sQ6+2G+5i5RKbHn1YfCNZeo82
qd9dAii6glqqGGvStV4hN5TiHftVxXF7L/MCb6z7kk8F8LMUxYl51kj+DkbVJG1J
ZYF5UNEGqNTpD71mQMxbbQSu7DGykI+ITa1N4vAgFo54s9iu5psLwzgaj1kWBGgn
pNEtHh9nxN/hauSWSW33lJ3+45G5HntnZ8GWnXZjqqXLUWEJRaVGGthA6/DGKu60
i5UHJ8dTcuoWEvmCmAUbGOH2Bgbroy4SmUoimLeQPZfj/GLTg6OTgz3hQB16SbI2
KBRHbX6FJhWFrBdlgSSEgojpTWFUXtK73RrkOQJB/MrCjh0eCi5ByANWoQcZuyVk
oDJPy3kqp8p/iONYRdZtSBXop3NCVbJJAP4yHom6lnzwoi/03eja7ouurRMDCnT5
mROkiF864om7EAKT6z7GWl1/OPjrEBaBiqXvYd4PkHbPc9vPsxzSXsLxn8IOEPud
ujBx8SoEx16YjUEGxQNhSicOFKcwWjMbeUpA3fGPOTTkZl3FRWKWlIe9jx1Js8dl
FaCEVnj1gWjpbfC4DRSQ8ha1ONVLPSUSVogQTRiXUdmOoCBPJqo/5LmArEIVsnsR
1Wx0w9xoDTbvxED574nSBdE2FjzuG0Z/PjuH/0mC89PZLrxLTy+FyTqy09noilQv
yVh80GkRpLjXYyaB8l0jP7ExmvzFloPaoIzLCGsXEW6bAhnaz2SJBKLOESGSrDo/
X5MYNDVF7WJPE2gxy+DUoMhBsumZZG/xArC7Qp20vaQA/Fna891LmiZdddmqC8dl
AhkbJ7NxE+xMpArDCGgq7pl1UTIvM98gWu470MopK2U9NfTD2evZAZh7Wd3kxGEE
kHf2eaj/Jcet+vF6/nUzHcZ+xE3ZZcDtC6QWX7GaddlDaV6tAFu0Cfb9M0Ds+rrY
EY3Fi3GArTQ3EwH5FNeINcPQaGeUcuL6Ylt38xxbbdBi5Zz/Zu3yk6dkkOf/r+mK
IEeGNBHaU5ZbUSdB74pgLQkiPaeDT55e7SjZV8xfUZIbWNeqQiBRlTCW3rlSKW4B
fnEyC+8CvUyI+yfaV3k5/6YbDHIz/BaILwOaREM+V7C8kzy8smi/0IQe3WekcTKV
0WeObkU8G0naS6rl9SjJ8J6+Y5WlI3o1HJTquc3b5iEhYqMZ4vCsAKLJoDHAE570
s8kra7NWKxYxWvtLftcDivBY+dIbslbyOfaTHTQd98l+zw42lF1FM3Jsfdadvb0K
mj5/NJ27WkaRYryQAPvrA+kqnrGnwj7HwriCXsk8nOoLbP2DjRCuibDma7UwU5/f
1DZFceSaU72jQ27GMx+J9vib1vOCuCtuVGjEZGoPsPiQ1upJXcSm04OPZdsocDs3
EttcS4xeDsq89JqdWQAH9NIFVohfgO6o6DbAIGkbaPuvp/lnYK8axML0LcAHsIdr
eolQKNUPCHL5IZjbVgfYtZLa7iq1Kx18+C8/QncVc4a4bYKUoNYchAxxy/WiuszM
9MZfdnB1qiaei68wMpo0ijP0rfRqc4fc+z/9CXnYyg4u0xwn9gSGsPDdjO1tdHVc
jreMmoyzb65zJFlFOY4l9V+b2/4BlZ6RUm3LbGi+ZFiSMj0S8iMccBFBP5fo93Wl
hHQ+1ZOmpjzAKYDt1HvypbB6yqhgqfy/wZLpQVw/rI9bOuY+ykyDVlCBlkIryUmW
QalWdll3WNE9ehZjHuF355aTvOC20GJfwOavPyMZj623IIKwVlbt5tm3TB3+oecW
om8mqOFT4glnrULIlXr+hZl5Gjhn9Q+VXSY1ilmTcrilxfzemS/y44ICLuSy9nlv
+slfizF4Zi6iYt+u5qHyJ66gRy9ggPnq2VTvwjODe/R7XRTSWKBX0AkviZsMTDEN
Z296SlX8ZkMMEc66MkgSBFgfLr7/ZnLZ67n+3JHuY1KnlyYXZfPkJgvuns0rvTOS
ZbSJcGFYWuxsbiBbgojLQRktN9ZDMMdDFUVvv5QjMO1KjvoHHYofscNXxUFIHUzs
DO3VwXBYeFUB1QyiEye6xA2wjwKSOy3NDxf8KPldoDMpvuTaKLRIW+yP5gSvMv2o
SeCtnno9zyIGmW+14S7/QuXDIo7OhNTIUpT0pSPUKPmVegpy2Dg2uTa/snUHb/Pn
pSCJFZlsINwerJTNbpHumSxbMAjdBkVEcWX6XvIWCHpg4q7i1tt79Y7ub4sHFQij
IheCdtplTQmekZEOgKAd6MuCUwtmlosIAVqdMfjA3Jh05bGSos2uS78AizEFwrah
yMwBv5YumO/q7eR7U6IdsngLZnI8vJn0IgDY0lQMvLtIFmNph5vrLdoczg3ro1l9
RnsJjJL7l1vqtDqDwj3QIezC0ar22BZvjXN/Kojg/0Eh6qW1vhYu2KTRn2hIrmDP
USyXoYq5YGz59POxwsDy0ZcS2Q2bQ34psCgi0XxvYPAnoHDqqow/OUdz2+R/7UJl
133TqSuikdFxkfI8Bt7HC16plEUYl9LEJyu2EweMQb3SEGSD0ZBPzpbhQvb9i4U1
IAAafR698GQQ3n1EyT9dFyyOnzCNb3GkoGtb7bSWq+uBxrkcaQsN9jYS7NvicM7S
ybHisvZ4E191exGfVKaW4dXq8DKRJ1h5otvBzZzDg00nOvSs0uTBPGA159Ud3MoM
lIlqv7y6eLZaXaDVDJYSeXAb0YRyKLrEP4q7DdhUJCQmYQmq9pjPZz2EXbgJE0v7
kuO32VBOkKgBa2k4L8KW+eSjOt+gHo1JQOneFKNcz2wxLGHKus7rd4EXTWAFj973
DE1MFDLMTTuSehuzPa/jfDSGlRJtte03wARGtNmRLoG9UZLxlOh78QLzJYpPkeGE
oxL/ET4TuAfYTXH95ILkOaaS/gVnjh8tY7ysqDW60Dm2/FZaFol6s7Hg2THPApbu
5aEAcQwYBG8cmAe5Ayf0tSstFbUxpqMCL22JzKeEUl0syYyPYZx60/05kn3z+n7Z
KkZNkjPwmMYFpNprYFK07cAAPwIzx/oMx4ynypP0AyVXNJB5z/acXLnkcB74gndF
dTjtCNJQqSrw+dvpZ0cELICokhNZoB+4Eq3rG5fu+7M9IA09RT8jUK2ZzPiJdJ4S
UFSwXE5D+rFS4LzUhPnxnqlDKGCNTqcJ9ky5e1Gzc++5g/Oh01CRORIxCJCqr9lZ
EcCwwjjaOhxg5UCud1m1fKvwEQpF3mT1Hlf8Wqkg5heDt6WZyUqn3/oI7hNNCDIS
2yap4aMhK6fpf3DRafakYQRcnBTWxsAkb6HA5ekLjetrYKS8r0qZFwYMFxRb0F1J
6kX+isSoATIMA7NQ1L87CldwRSxLiqeRGtvqXG4PBDwFaEm5d9GWAvROW1v17/b8
jwlq0HUeIfaI7E9oK5TUojIVTFWnFB+0g4Ce3Tbt7KgCXEgdfyKoV/7W/O/UTCY/
aJmjM+PqdM6PHgcDEtBkfZr4KLGuATjzeWSBy8u2L+ap8wlTC1dWdNQAAV/AsNai
8nkRXouWq10oWNXu8dzyz6YIBzhcetdpGRzJmG9qy9PhWfHM780wAPFkLyfdKOYH
HoOBToBqXr1PAumsQa2qL0xY8P26zx4WA4isdpytpmwpqOQf2EFbG4zNknfoFEr1
m8DzD8NPB/P5LqXcCcQx0CqFA4/JnvKGZ6SOWBeI6789br4axyDoco3Qe8/GZON2
U4hXzSZ2dKgZQt/DyKfgohFyNUjMuS3daHZJ5BVXw/LfibQszVJRqhzBQxQVbYDl
F7EZWeSS5CZAH5gtZGzLpnKKqPvQ2v5Z+DKDscj75gaHk2uOMO71EEiCdx5KOsG4
kvlT5yxLQmZ5msh9PEoH45rLeOOEe4dgLUCD/rwdiw/Fz8HGAUIJsz8N0G3uA1lt
Q3qrAPwsE4p8Sk1XtuNZYaaq7ePO6TZWQ0scz4yskhCYenOW916BU0PUmTNAn78M
G+zD9uYo52iMvvEmufyYHisRw7LVTVGYbUAU5WvYsvEgsGH7XSmsERPxLQBColWm
lVCYADU8qZ3TxRucXtlri7fC2LN/3FyILHsY2oH/5+UBQ2sWIPdfHNLG6s1RhrTe
mPhUVKlnv8OEyD0ESdG9dH+VrksyA0SEoOrypsP80U3tEpSEX40OeHq1lgNBZW5J
xQLZBs80Hmnu3jCm5KVALijKCXPvG2uUH7G3ds/DYnOSLiT7AekTdQNQ0v/fX9Xy
TIQbvWtfHB+8/4wH9V5qpCRC7qO6lrRbJM5oej2sUqRDt8qYhL4cZyV5gF3H5drU
MknwhEnzq9QryHijoVcRc3wENACtm48Gahctys09S3adJyyIIKaQfJBT4EEik8jU
dHc31IM/AhPFdxRZ3L0Hf64Zd/841bXFKtVQfkVZWt+wPfAQ9IBNoCC4Pd/NJ4dc
XNhLLgAn/oLDRxagKDHEaNAuX08M/cU2zaNtdT/+U2qExtDH+7XPZgGCnsL1kzn6
HRUx24v6jrEC9T9obM+inZbG5su2p8csdHNt2slX1TTUNfZ8IGOICB/OpGh1nBAU
OJa/71qDHHYIZ0wMC9TQKYoeEHB7JhXwiVF8fVVWFjKXzmXiPLEtNFbZ/cEag8AU
zsYWkhnIPMlZBvz9oWmYXpwaOzexXpdqNVJygKLdU/ddURdNYGV8R5G9Ey14EZwZ
9693iUxBM3Q/gOVuZAOMNBR+6GpLSpxDunJmo1cGX8bvMDf9VxwdWQ43tstwCEEr
lAJEAAP/nrFuBcdZ9D75ru6AAwwl62rwEhgvKbHjFbEsMQVuEr4jb4cW9ACL86ki
uOrajjssnf11YMwBLBMcmUl2/LFU526Ht66zLd1VwvN+wFwKQM0sOS2VtS9BQet8
paTPNqxbEczL2ecyGuQsV//iv7DQe3OzA2PX9zFEoqqLBQjrJpMrW/8u6HGEka+D
bWdbr/MLYjWCGaeFhyCYKjc2wroUchfFO0YHBfiXQ3JtuLjuix3Rhsz/908eFMpA
Iop7Hp0hgbYq6uaA38ijkagxcYNWBb6L1rbJBcnoT8uFHGGSh3U2TGf0UpEkhIsz
AJ6YIIBD2XDZMaVJBUGtHA0vl1ZZ1BM1MTyV6QVovKmyydQz48YXnPHaGBRMikQ2
UZi2W9elEfDaWUk4ULSwZATGlOqtuYxz/dhWd+zhiLb5y4zBDG4J7aBdvNxFbFMl
ImigNC4fqrL+HfsGIBmDIKPpV2OQlnNj8srFqY7HN0JolXTRNlc6JtHOb1Cr4FvG
3O0A8LNXIRYCc76IhDA/eZSvRcdHu6AwAe/v2uN3gF5AQzsa3bHhYKN3MIMwPCA+
SWsPNGw6A+qjQLfXuvG0HgTxMgn9ZZYtHMRWT4F8lGXSlIcNZqDmmQWgzisMO0Es
n70+TGok9qE6H8/KWgMu7Z+AesXf+WqxmBk11yo+njag3lfu/XA27/fdMKJW/ceC
Finiop6FGwwhb8AXoH2WWs++pRAp5ml7AbibpX1D83eEtMhFiGbHii40WhMdcDAV
0DedJqB1rsnPtqy1HOghdhe2sQhUQ8IcaimKVt+XepJ+lvFvDMoR80uGmz69NN1E
DvPWvwakIu/GtqoqZbaNZISKKoFW2YSVQ7ypViYDWV/YiSQtegLo55Mrd2vUCCw1
qRHYVwCYBb55QSKvgU6lkP/Ay48hQ63PKHLu/z75GFZaTAaf3tMtEHy8LqYlhONf
C0jy2nidSErHOz3UWfNMcAzw014RWGcCKsAn/xgsovOrAiHRH8vH9A49G9bLjysj
41b1Fe9a62G8kosB6R26Nc3FCk0Lh1tYeSTs3OmfYodO9Vg5ifDTgLkOA35kCoxG
Ub3bIQu7DTZLYeiu8nCeo4KCXde5MTn4k0Vf8kn4MDTF4u4af/H0k7aBXTSF1JQw
6N9W+y2VqDZiq6eBovWhHh7EEI5+Od5m6nsnydxa5rUGD01yy1sfoiw9iXtd5RV3
INwc2qOfGSc2AaZHhXq09ULnihIaAdFTPj9QxFHSTnbdHPZkaNNeyIgT867Hwpxi
XkhWuqDeJZjNQN/U/mK/nKIFoRhNfvXiHgkoe+eYqM3y8k7kmUDQQ5LT3MlUseRp
KuJV5SNddIUOyKMy/S+zrK6LT+7I7zzz1Bg7sH9/SwlhpQgiFuiq3eB1SVqZUEKR
coJjxShGnSTTV/YbKzhf9XoB/w0swo/Cy9MpcSFR/i247qI/JQIPd/8TGJW/hrnp
d0bQUTIRrIBV8f0iF4Dv1tO3JKMPUv0PjEWGRB+pmTEha6yUUvz0lUACP5pO4Ygl
7FR0QiAOXmTXua5a7H1CNTdoinLmm+BLHDbZzsaMMKS68ib6f0JrQg5HdWVBa/1B
uvtYNlJvqCaLc7z0KQ+z8GN8pElse5fNrQYH4ETGEUfB40+ok3alOhQI5roESCDR
TSTPslNNkX/YTiFTkxFgzdEjWEE5l5xHZ/qRBw4JiS89W9p9+d1M8Yv6pS5d0Fyy
M7Da/DQ7d9rCZ+vyA0x6qvgzz+qklRT4Y4OC9FlsB0MAEhjk5S/J4V94rDSAFMgI
lDe7MyCjT+z/Ym1apnzu/II/Hd+ILJy6UH8hY/3EZxC7c/ORJgc7HjjrN9f2iWmF
Qdouibm+N4+w57wA4JpXzOcuPJLjCYTFyMmAkBV0Ytr0fY/qjKC9nycIXVX6MUbB
mud+nQh22lp9dn0yv3AY81QAKDMT4XjXbgOZpTVoU0wrAXPB1wWsm3+e4904TeAN
gBrVAFiiVvcMj5UgwxCkDc4VyLhA794+4uZJXk3+5jUTmCaMNFeizdmokQh4pM8j
cZOgbW2320nWSCeLziG8xA8C4HkkO5g/TFTikWAp4ovmwj525CwQpQMEFwxeS+Rt
gD4fcjZ1A3RIuNlO6PJ+QkePpEW//hkMr9fOhcMhOW0YIbOBsDPxbgv+h7p08hZT
2RcJzKPWBNkOTRzS+mGX9k0nGB/qZ9HX+4FgI2dFZcozeoC2q8Hv6c0YQGCDKojf
+GwgaBEsHKPUbGp0YNS1wi2ijo5V3ikm5kC7LTdirRR/nDfhkkiEEbNmndiuzHy3
7RCsk1eyLD4gEKJbNt6oRhJeo0uHyWNijD4FgISKK6KFv5EqAPh2jAVJQsgRKPSH
cbR48ghfTeHDrkap4i6CzutEMfgBwkYLwUuTARJSFVxZLa/bOWG7CYp7sS8Qzl7A
LKGAeKM6O4S+ZTgSHhyIgaoihdhxNKEMjSs+Wy73/Ha5Q+itniN8Cs/Fj+b5TFSq
M+hVmbIcvGaE+wFGrMjhUjli6yQxPpfdeGkd5B7Juma+CQ2r2IMO2eRrwQdYAYqy
oehXXE6HTCoBzH/PVdCDY1SqoklekWQMoNQua6ZmE6HkwJiDtOj5TiP379jGTeBu
JcRNQw05yVBqC+2WqFm+B04dxRXy2HdzLM1skhvvjCds399HICXnHPXXiWgTD/1Z
tHTDPcOq17OwnMs4YuxBPhivJHxAC+s6joMuTG3FpAv4dDrPXkZG6GFpwQamB7Sz
ByIiCpRKfY+x8fVfN3s/dCRel8lmt6tokIgjU23RBKvUB5NAjw3Nrrm9iKHuEsTk
TvDqmKoiSxj66pCPo9AdErh9oCJLjSTEuyd9CRPCoqVtk8Yb/lF6oooBaSnxIPXp
fhw0Qv/y1B0FTUW3xF/wLmRWi++vxOa/Tp3Z7YgVQhl42rLBfddRUfXDagCo4deQ
z46Ru2KAsyJ1PIX6VKKD7EzL7PQ1VLWyyobfagwFfsTFqmuofxpW7gJQlrgrI0hT
p1vTnkGWBvT9r57e4V16cG1g8BVUwZniOPFudtVvhG8GTZLbVBLqB2MdSsE3lt+L
UkqlETFRlLaOq8NjhJbFoQ/7O4nJEmURRZWG/kHnQhhyBXy9QdhUYgORUpUKnA7w
6BnzZvrcdpETenP8wOB6ovhMg0gmUGMsjTibaPD34g2c8bdT/p2ap4kP5xEYbK0K
mWTxjkqpSLSVRtLX+6RzCvNomEZrWE8DG7/wWZK/zsdAYjtBYzaRteoMJoVuuZo+
zo3Kk6obUPZzmp/lM/4S10kNbNqoTiDNTQt4VE8TWL7xO44cyzKpbb3QOw2IZRtw
Za9MRJgXZQMfYwhlMCJM5r4qfVAZlbrMtR/ZP6el4y0JqdfB7ANAg3G9tUWQrs1Y
4mlByzIMi1Czz3eK5t8ubvpQDFWwX/IH85F9oADKH2B5CcxCfgV6b8dqAB2cL2pH
dPB3hn44zwTIou838FColc8/Jvg/c50sLqO8qvHl4jNgDaOpoJYcqlrWUd9DTBPT
MMenbn4lCZQUIfE8NU2iLacwRH5lT7zKrT6fW1TMC+ecTZ4iyEaox6uz5jyziF99
kIzfWda/yyUUuyBkh3wQWKHLjJR2ple7s2jsoOd0pavLjC4TYWdSpA45DOLa/qRl
kqYba9pYDHpFYlG17cyU39FDE0XVyHufCIlCexSvMYNQ85UYPrLcn5YBerKBP0RQ
RaMrjaAFw9tFhCmeCNCSR60Jh0QMMoeq3jRl0OC6EqYZOnfkD7+TBIPLfOYSB4b+
IfpPraTlkjNjCAD4wnOWUq5IxTaOboh/4fm0aZaGYnpcS3+x4M3D+8WoBA5ZLSmL
XzCFMxNM3I0kPdwF8YurdBO0Rz/aYQ1yssm9IkENh4cuoX4+5GBR5C8rbU0uR2fY
LOvOpOWCtONO2iaC7UhumATBvM0Z4OhJwDGVGVJxeobMiDP5/YG/b7gIgxk2ljbT
3xN5iTOSwQfIVb7c3bNYmzk26oW+CXYD7PJhJNM13OoKoF/8jwh4HZ0tGCzSBymv
NrwdA8k0fEZ8CHOatBQDB7YilqQFOrIo9wTbiFU/2sxyxL8+c4Ni9+xhdMtpoA2K
kVu676scgY+lRTeYzl9wshxk7/vzkiuSMUYUtEjh8dmGJDCWX8QDa74DZ4tlOoDQ
WVG5yB7LIC00BXt+9DppdZlYbxV7MuzWvj5vU288RZPBhPd6MvaFPoqkksYTfl5w
j7lYJ7m51FFrRt3asKSx29ogqsRSsOGiuPuFNnFf5WL+loUX4aageLQK7t9CKDPT
HGU7vgLs8WTQZ9rG1iNhtaFyV1eWidfGrk8Hm4wz+34dBLmg8H5abKmUKLxNqmO4
z5LBTTuDkd3Q+RDWvm2zWSbI8EbJ8ZMtZAx+a4I+/oCYrXLfvmmvzUBzpXPybVQ8
hETVTxRCEChCg7ZXSHQO/AGQS/c6WHpHNSPaOQbQNPcJgppGtGDFfL/XslbOIh+f
uXmmJLmUkPTxl1o84QZV4A1weMmfkOSIcgvYYfkt5fzTkjrwZapLnxLBBHOP4Hzg
BVrR+/JVoRCxQpt9V1s4JOFYZG13vOPW1XCwTEsADxUG3EJKpxhny5hQXGq8zsiQ
NKp5L1wT7JEtjfkMGBasEu1fHVcx64oNNo3s1OofUOXwyQWoC5YBAgBeFLsaLBys
DOOBY4LFtWnrudRQ6qipSuGDghqKx9/46kPLdn7hLyGy2ml0+9JVtm+GKEvZfqFS
ompnIs2Nb9lEgQpecipWkEw3jhJ4pRNW4R+IzZYC/G586CNdbIGHi1Khg/+si7re
uho1xpq5A7sBeN8Jv2skzXA/DRN8eL2mTZ9slm5XvWkakSN/66LeYPbG6FCs2iw0
19ShgXQ0gio4ILdKsgfve0dRlrd5FHxPC9emhOVRin6VCEACwwfyBUXKGkM9CEuM
CtjkDC8EhC2cthy+BKHeI6f4aBQCx/hRLyFPgMiYZak7UuIgoYoY/rCTTssjvt4k
zyLzpQP+AvH5ktrJ5zMRPYc99WmPo+WhZtFAiqgXGHhT9jIatPYhL2jHMC7aEDIk
DkMyUamObM73vzqrL2Kw11fy9+hBWAltW9DNy7zoyXHUQfvWosO9n4X6HtY0j6HF
lyod9U5FhtQ6KrJ5fi7aq/3tjAZQK7ZeFk9YP0QO/QunveGlFJe0c0Ydnqlgsrrf
FvVxBgnZTW3sQjZTnMJ0yN1gI8qaQPPYwn2VzxrxC5hzw8jke8OBVdY/FDDheMxV
B+ZD2RmulLbTh8jFYw1S7hHTVgHRgTyuGeYA/xOxU6CYLJy6t7q6E11Ai/E5iCZc
EFwFOC2je6zLPkanMKjG4tfsjWZ8iJWIPyxMbXuqQNZZ2rUdbnSkck2IYzt9jKtZ
UfOZHUTmayv4yS86mPOgVl+8+boJBVRXE2Xz59TMw8DVkGh0/h6kr03PlzBzJIpG
vGQbW+b4PSOYHTX9ovR/aINKKm5c6Sru8fGjxU2z2zZK0HR7vWKigv5C9/79MqZ6
Ph+KHsjisugzrFVQ1VVmsFLJW/xAzMZebRgHcrkM9XAuknrDXz+hd19RHlAnL0cf
7mC8vhJvYrgxrEdg66kAgg+94y4Oc0+catRVEHijXKJOjVGfUGgG3QHC2ychPhiQ
cltxaenHxV9fYiCMS7cvlhiCM6/VSSHmdnmYF7Ojw6gp7mL3QeI4Y7fG4zsFiI1S
o7z+JHTZ/OkuGasBwlhur8eFYmCQvE+AEQiu0k6HaBuq8QS3E2khcBCy6DiuZN6P
Bf7oexGBag48kI6rGortS1uQxfCuKS6CYfhDoFUqHxnLHE0lun1v1fGwqsxCLYMG
Dm0tk+vPtczQHC4ul2G0Y7e45YYB+CElCAQD5Jv63rtCngpuJm2JWfA6G4SZPC5b
V66u6kwUP01m2ZnvtEFap4zMjOGSP2Gi95WEk+qzezcBlJrEuTh3AGWxTkN1MYUB
R9CJ9KmhGOQ57k+EFhN+S/RKS7M6SjyZlU3Gs6bUtrWq0J8rdfYuoyZ8qfd9D8j7
hcIP3RO9aWMxJPcHYLXC2NHYuYBpjHFIV/4b61Ik6X4f1ZCbeWqWTH9sEb+Tp/hg
3Uqjzo7ovp7iN0ympSwbvvQLyvOJtBQf4eAV89MomIXJvUVr+5MNgdohTrpFOLiZ
oq3BVaRvGs7DZuflyVW6l9al5P/ArmMy2J+aU6Ljg8VQxAtmgf3ArFuc60AHMsnj
U+V042Ja5Mld10+StG7l4ETubx4uTqtOVQru1esU7BVDJqwmV12SRSjKkH6LKtZv
R0zhrFRByzKyKUm1rOtVBCB8id4HTzpjRnCUYqPJ00dlpjHmTutywSiDgQV+kEEy
m3Jn82hUAVjvwBGNQEiXWoZB4Ww+cJHE70H/LOynE9aVkX7XyrooUdwU7RgpkCOI
G2vIRIi/mSS0e3tCcrsfzjCBZvTwCATjqUbcyIIS22nnnIVPSefjkACVQuGKo904
dbmF0kJDawlDWAOUegEu3algIK7MLpH7sdklya065hUpf6lbHxLaqPawp8E9/6QT
JuaqADCJRfX+DVOdzpZ4oML5ZxQLfwSQcZASdQ1lKLz5rOWfRNcWLat/KeXxZfRq
Qo8l4Xtx3E03t1iSA+5qQQZ+R4CSiQ9N1F6t5qsU9H/PiZlV6MOvvCgWHHQapzGm
naJebuzlwkwlu73wwUwffHWLdtx00Ib7E6EXzoc1HQnYjCn3ZPWy+cf3O38+iQ3i
dZYBZlVD9FmFEFydWGQ/Ujbev/ZZ/05qVDN3D4ce/m6iwclICSwSdlFi2e7J9VR9
4vIOvN758JstrGdwOlAbZV6/VTm2rR0APyAiz0A+Tpx2IfEqc/JcL54EVYsxT3xv
5N8xvlT9utyz7AHHr0vBjOPzbtGcAswFWhrra26Ec4oPyrPkJOzgxVkJxBizvSen
jtwgxdj6ZdPjsKlqSlyVcgipDgbUA+XT9mnhNdeHpwAt81aXGAtkO594BPniwCuH
AT+pEzfjx0v3pheRtK0q9R89B0X7cdY15X+PRQuXWs3AUJOsDkTJbQCfLFMQ2LfA
gLcML6vZaCf8PVrYvbobUk3V1JXteK62x9+7Opq0jlb0EFq9VHvilhv5D9WcO8Sb
l2cSLqehKufyvx4IDCtMX6kyKAsYnWmh2Uf13+iQQ5BncbS1AjmNEL6K0Z2417rn
0CLe+bZLNq+S4zUDf2IZeIuGqE+bMWl3mL+b+vrFfRLxZGDTI5blWi5lXCDyeddE
hGuDAD8VNyBphrG0Eq3QOYXV/a4GeBb7+UfVk7LPGaI8+tvUx8mkGmd/lCiFVTWV
/In5/ThM9E3FSjfh9VhzL+eAFGs9aZ9HZrrT52WifCYmv9Ovb2LxCNd5gTDu+N4Q
Tkr2ozqzc+gBnrIfjOR/Z7btfs4KT6mTeIeyJCCvlTqdsDC6fP2wmHY4CTBlJ4lc
0KMF22XPNSHlOn0tt9rHiFt35ulFP9Vn8QSvNYWcpeZUwZM6euU8eYij+eGHDb30
jdcs8hdEW5cFjrXqwWlJjO9n++BkQMipvRREmrzha1zlmYPchff4lHgzqCS5ZYo2
+mSXdSkH3qok8otetEb4/2kbPvvjA0LWsPCLjXGHbz1jMRjwfqKIiDi4nJIgwoIG
GQ36VPfzTvf56gtenubmEGSMEJer3k6Dyf+jSxlYfLhL9HpAyew4S5jb18LfOz3k
6i9F7w4CQj8M8jOD9Wsb6tSAcUvbX5H5aBf98DzX0a4mq457If51USZzp2wNfreI
rUMkdFLoX0Q75iEz7sDy111trY3vCEQS2eF5b4b2KVtq7jANOehXzhqCMBgh/06c
Kh+GX62cGLly7npEVJ57rzfx8L0cr8vCDdck0A+PkINzFOcbbG0WrtgI8eR1veym
/0PD6tF3RK7XD09v7qf0ltlPHMwVh7qfOYtu+QAG8BXdw1QPDGxXCYfc6at8vneq
pgPS8spzRgTUuQxpTJIYVRmsFEYFgm951FyCR/UxQ6lq3sOvXp1OGA1kSzDAozNV
OrpwNWzQjkrerNukvY55V1qDDuq7UTYdY+EKiU4jBgNSsh5xveddpzg/zGp+onDM
A9UBPXc46DtmQhFs0wsigh1Ig/W/18GyifyxHq2fO0uucC3CYw34XYIiMjx6AAug
Uft/gouuqlkj7vO9768qdYcg0Zk46I+TrBWHfMYdqnVtAANU74PX6mH/ToRXvNB2
4GPF95YVnJV+6qD3F78euIAYNExjnLRvtMJhhCZLLwGsDHT2yEbHIZssGjhh8Yir
10f8c9pH3bb9irti98fDYhwyxBqTD55ywvPDVY4tsmxxLW51R4RDTgW4cw50wKkR
uymOLwT0M6zNAFR2wjUVTyQayOL8Q18azE8W1WAcGRf0Lg5bsPYtX0UWZXuNVnyD
1/mpDHKFupx2qIS0z462xuhwZ8/7/wV6HK8FuoAjLwBfc1ipgmIAJlpdQ4ZEt+nN
ef2dF1FFAp7GWJlk4L6ZtMo/iduJJdBf1B0ISuvZZ1i96va6I7zwzmUeVyjP6DQY
zX9dSyHsLUTnzFdzJsv9guZmo1RLGTIm+3qVt6ZIZRdE3TR2FvnrQnv/qK9thtur
PXXgzN37BZFSn8uKELQmjCbPsNhfSOx7fLi6Pgm53WlPIKhkeF1OhS2L8O4l0olu
Wb03rsgWL+s5r2YmDTArrdDDBLgSwnRpk4PES2XP1k4LcfGWhnoNV0eOUo9WGgb6
ya5eBy6124RFUaFZy74sMFwT7I8IB5ZnHd/aKSglwqTkZtH05cyr5JM71u4KMRIr
iih29fTnDtaUyaMdRPlSqRIHV397189qKtec/kxNRFpctbJFgpK7o+wj52GslEWb
rnfr0/TAvTmkLYT0t78/S69ONlVsXziSsn7P4TXv2oS7sXnNZKB6Es5WGBFKRTbk
tnWqn85p7riY/pw5qxIJe0sOopvGuD00fKBd9LD0JRwdWPt4kwGFS2/G19L5f0kP
bJ+Eyyrl7peBhqtadt3R4hzP7bsvnPrm28taUrLX8j+p8RM8u3uF6O/uxr/YY/zG
h8yTLQfpT8kvJrU6tCsPkzaZZ5Ebu85D7yXHQt78Cnq3Vd5SzFQ+bYiMl2zea5jd
5M2bXGyZn0ncVnjQ+xGtvWHbkEorV0FEasbBhckxOM932Cp75twkFe435g6+Mgs/
oSRag/RwAgLA6M+1hh1wAyf9kdxsa4LUfymRq7GXe5McXgcPqJ0QArqCh9uiRfL0
j/yVMKQ0Yp9I/YPMvcnfvGFyWAGDWoL9KYNT3UdZkHnghhobkkRRwoJh+ygRR9iV
MpySP9EHXdxK7N9LWGyBk4Jl56wNeJNhN5cbI0qQBqUH7OQ8ydyhhTRZCzPYu6GN
ZcPRgHB0U6G5Qsj7yhSa7U7tnimx8GYSHWBVDVCVm1K/WxicQ5G1trAHw93ltP/V
S9k4cPTR/T4bavPyNC/swfXdjvbak22saZO+1NyfBFpTrfKrT3kSnt1HO18La0jF
HWXB7q5OWGYdHVYdfqiGvJCGkWVxIgFIdded9n6bCjMWRfAiJocnNuoC8koWPRuZ
mHU4WjiZv/qTL3Hw6g4joKdIdI5QA1FSPaB7rHLcm9SHsM8nsa8KEe2nQ4sRg1og
4e5W1stmN93PyppqqJc0YHNvCOnL0T12wO0ClU3ooV6b4ecViiLyuzowchwfmoJI
1Not+12RawtlldrObiWuOTlExEq9J5zfMHcO0PXmdqCtZpDxTv/7T9SXsCXrzm8D
VS3PG1pDPk0awmG33//ksgsN9ffk69zIE3T1rd1X+Q5bz9/BO0FdjMhsZo5T+XyF
0OWXgay6R4bsoPhMpf8Efzv/VlY9XztFrILZ8lLtuO/STVcsfOHR2B8FEitNj+uw
V3sspe7lKWNB+PXtWinxe7XP9EPRGL+HQ0xYcifUY5tQ8L7b9aIwiuDDzY3sdFkM
dTonKPhI/KIr0/VvwW/DsMyoN+ATHdoCbS20TlGjWgrGXqVQsKH5ahTQcDidkrGy
bYBh9ZN6rtDaUchezl55qwTPAZEInsWho1j0v20xfSy+gQvj9KqyhV8y+lHbSVno
xky9jyt2zf3nwUc2Mo/UsWCpYj0wG9L8CaUaFGRyHtrrZ2c3O0ame4hoRXZTavg5
XF5w1QrCkbl95SJ/ItR0ntKoaT8tlGi0H/0mYB0zMc5b2UxuxK6x+PQC9pvkI645
Yys5hw43qC/xG3gYRfJmTgOdV9evtfD/AMaP3W+NIwMjYBKBdXNoUrczUyADqfVO
Mf3gFO/YsuxRNUa2+F6p+Kbw0HnHNeE4dAgNco9C2jf8jnFeMfshfr7r3L4HVkyx
zNicyMA6s9iOSABLs3+wFQP3n2tU8SnqgYkY87NMKb9W6Q+Qqi+zOA7J27Hz1oij
JwWGOfthdQ2XPbuqhv0yx0MJYcEkKgx81s2KDUyBwmnHta4M5vltUCnGB4JHgteX
xysNzA1mYLYiWWr6z388CB0aJFzGb9GYmVuJKTrGvdbS2MSZAOcPbLasGIOiboGE
jWIYRHMvpZNvZ87sBO29YPQk6XIPnFjRnWfu7QjQ2xXuSkz9kkaoo3TxQ2Oae8V2
HyzZOaykMrQ0WO+aaxnG3XRLbI5wex4TSnOXl7/EZUHMonUWuQzguNBfWtbusda8
UiqGPfAYETHWm7vdMbe73DXaOIsCMrbjZALOzthinAtUbiQ+aG0wUiSO0vj1SHF8
uB8gY0oI5XDKzeNbmfuEayuCuNdKp20hfxK+huQmpogLpkfYCb2ksHWqNtYJyYR8
fSb9/17Ce7hw4oi7O/mKW6r5MTbgwsCIWZ9phRS7CA1/EdxMiXZ8tmYcoKWiVxc/
7EDY8xgU/YJsDIyzAYYu55rZvXMtiuz1vZ157vB1aYzyJLZNjjFBBck67n6LuTFv
7Bf74HgbriePG7zl0cmn1ELHMuQPkS5PH9aieu2DwzaIKqHLM5bgOpoMvisGk6N8
ac+xZCcGaNlqBpJ1Y+1ximuZMmAqqzBgw3nOhwm9JBoMjbRaxPLXlBndHEzxs+2X
1Z0npMeq/lCMtF+BFwnfMYuS53awn/ueX+/Yb+GJm517zlehqLIfYMAeno8Wn40z
0itds0+b40O18/Gr/duTfpzMrWDTqS5dc4hHjCzTlf1PXYRSyathH5LzN2UbH/fU
h8FVl60WNgZIOnA++zf55vfyaY2ilRTrvhm1inPrfBFOUrOy8MUNtaXPpiHWJzhk
JlyrO0RQH4VAN+BS9VP+G9+eLyGF2ScozLizLT1BegOOUSkqPWQh0TWeeQxF7mSw
8jV12ptePrVOtlJZOuM1sM8MGS28BEUF8NBP7WAHmvqvnjDmFvv/rUpP8VlrSPpx
1PFPcUNNVAcOnTLRUJA24MQUoLVBwCKK6mxJtJpe1j238X6snlrPks4nHtQCzo5W
XzC310awS9dTYXtFaRCMH8VPJG8SE7QAIsGI1m/H9Yl8S1zBw6gZf1QRnETzjPkH
DqPMvKqUbNU9uad0ZcdLbiNXkU89XNKO/475qfMrxo/bDc0sV1o54FkkFQjF62sz
4h/80huNHkYM9q4TJMSeMcPLajI7NMukIMgcZU+t9Lk0795bjgoVJPg+qqEbwq3Y
wARJkraN9limRx+pXZyVrIxRsUVJ5ROlfC5rknThcidPYR7YlGvEcn1QRHmvakIZ
utFBYwws4BJPSG7Cr2S+8Qx5uxPhInBpL3ghIY0zKtVutzNr5xdExomD/OYivq0f
iOY4uUmRpCoWMr52p1SSKIjnrkIwsCz8zq+jc6J9nUbxw3RKO7DwbZ+WkepHuovI
ph1AWOJPLVNgtLAIQl7wKpXFqHL+ajC2LnDTZow6DupmS1ORLscp4/zkIe4ZD4qA
ys2xBuo4CF8p8+eyTZKRloAa9gBggOkQxcpCV+7WvSaZmxS1QxzngD4crp06p8fN
1g4ILNOD+9SQf1718JUSjaVtgaPhN6vCjVjxe7JXVkK7Nd6gF7JZhCGFi+wV5Njz
nThXSmKw1sVckZo6CQM2bBuP242nN0MF8FOpgxrz+dHEOcfEy15MyoxnNxU2+PQN
z+w/c4irb875OvmRcztKFH9YjZ0+FbY3FH00ValT2BtIloTUwiL3DqLlW5NvVm/n
Qp6ReQugmUtR/hgqiATWT8r+nFhwGwgTF46NV9QHIlDC6628GFS2tfM686WKDufg
qDcawm9FwQiGM6soTZqVaX5Tf+MCWig6MIJf66JzzwIQ8o69nK5RE+3e2XATeSGs
oli5MUJ0DrPEi6rTOi5B6AtEZ5Z1YHqh13JB3koWfpCMnbHzogge3I4V7pVNT0+J
vNxcfkHke8mLdFivq9h0QsqD5+PBw3e5NBkbIjzmGOY1OTQGL2CF/PiRgJN8mTA+
82WgaNj3hi8+u1BNtPlyuFWtvX0XpkVFoqYm8ctZk66tvJdWhPvDA0eHlxSqI4mA
s6My31cg5sectBR4i+GOMHSwvYv27+bVODaaJdOjznu62F21g4JbKkWCoH28Kss1
BXpu9b6JWB50jzpoV2Z8FMXrthCHsviiNdLYZ8JFDW1K75gz8w0su9XdRroymbMh
HLvwxfJAvmwgclKhfM0tocoDJtAophEbDWRU0XTPJvJE6mLVWav8aYuXuGzvPHSQ
iez1a9mFN0cZdmC2fZUzm5SBgPqG9NYEqEy0Q1WHqa5cEqbvjd0VqjS20AOaEKrR
DTCDURmwSF8Ur+OuxgP9wAumEfe1Xp5vabmrgiGS9WBMaNo9vuEJA3w8wqlMAMe8
+hOc6nlRvAdlHHH+QqZtKT9PMWFqGXFM9QYh091WzLTPpQxndNHxsmvGPIre7L04
FTW1Y9tVvfsP7jhmvbHhKFkoNhP5REF43cxwUg6zj0HqOThhyA9bWbu7tPm5g4Wg
JjLsvuj9xORTC3RmObulxNyxCkAvC6XJTewf5CyND9CyILXKbHKmUa0Q8mlMu6YD
eDWeql1DvnCgTixFznXAEoJMh2uEWCykNZygvqqcjAeXZ60mo3oWh6+Nc0H7Dn2F
gn8/aIVwDCFAdok/NHfk6JIr6VjIVrEWyP7ic5jsjEHjPfnZU4rdx6qprBiwY4br
/zIwahXK3nJTNrHok83bKohzuLAjTW2SyadeS3LC2yVwQUUkWE4UvdXMeB6Dp2Ml
bCq6j6oyiwmoei2rZsEYJzC26F1NaHAIPzVGlBUwkKTVt2UbH26I4fO0aLwTddcz
X5KP9tA9ImRXiyTg5haYp3JD3mvNdxc5qt0jHgJQtZeb6Io+OXEStHjSnOED4wpg
TZEFkE0Pe0mA5c3/KAUd98sdcAowiZrcB5Lq3Nt3WDjMf0jn7DVG4RJqMeC85YJH
VtyLeo07DA2C1SZBIeENqZlUJ1BxW0QnmL4Yz3e0uQcmo8MSbDjHErrCEtU5nqkt
zR8HuccT4A13EZm+aCK6brFiIsRp3UJgZPZX7EjyWtbpwA2G8y5xfa/VuGgSimNE
ypZIZSwK16XNdwQphS6LTzs7yd0oHMVAfrvl1QGkLchxWktJ/Xaba+xPj3t/nukQ
GYLT5hR80Il+jlOxw/jcNUU/kHbbqhEzXvp5fWYFRtPal3Ur5b6rBeUuuub3V6uQ
TMqqkf1an6DgNyGZ2VVwERbVyFYqehkRxcekcM+ge9vLXWswVbTeUUvmmwII3x86
KyiTe4dELnUE7yqfdnve0d6kbQTHkxiYH39O+M5wB6L+nTqwNC0FOqX3X29z3dHC
FXXaSt20v3SJHpFsm8lgU0QCNbB/89tiwFlELnBisxtG83jSTx6k/uo8kDkkh9Hn
YtCcFOq2TbJ4jpZU8npKqe+E1+ooN539OmNouugB+NBRd/Y180rp8g5wrXIttKyq
8eD5fDG0cxRH2Q7jzpfzSJOZWcRonL6nnVwE9mH6Li8IMRhjXNYRxHlWHONUHhhU
rmDs5DB5R1PJsMxOOLimGF5AUpZeBHou265zhU6bqHq26zwb3Lay1NtKjVuXoF6r
fKVdb7+vfRYl1C8DCvPhURrOIMceeWpECQhiBkawy0dZvFxtPKDa0rcl4+LPxVXy
morCQC1NQjRX65Ja+Z+qIupM9lbCAVR+SQtJQAC81UkGEyo7tBY5DxqZet/SljmJ
aLDlcaQ5nIoqy1CZh9WLxOCaGA/ub/48kYeEF/er4Pc0a/wC00appcpgrVDuAJNW
+PiK5OshylwypmusFr8DzKcyNBUzAp06WjK7p3oLYZomSBzlAk7c3UHLohrDSyNN
/JbCKWTljQmbnR+yhY7mzO0Cj/jVrWZr7YO8rCiEuN2lKsJq8q7m6ptL+kuiAF4t
vCwZgRFVQbtuEhTAaCqOnrR4D3dUa0dvYg3cRRL3Zv4dcpWcRoYavvgRxI5OCRcx
NLSiW3z9C7PGYmdgN0QUqlCnkZIRXP1VBKBsqz//EgDgRZsUa4WhgR52EbJROiQc
tXUl8H6vmfIq1mnY8wWklNrMDkJ4GCN09IZ/XiwknG76VRHYAtStCr945lDp1sxb
JVeHCmNo6MiT9dg7pNU9TFMOBmFCHna78puTaGm8m1FdXHFEdGCxZdSgaTvT087r
1ssiJM0IYkR2+FmCMfY9nuxTiY8u8Kewl557FKsAUbVF021ZnAHhmoWF81O97u2s
SHMZ2YcQs8l0G8NjkZ5mjzVxrg1g3i1yFpNmfNUpZUEbzxtLZQDX3eiIX2Hxk4FF
v34FW71ng0srQoqNr2EDzpoMyDoex+klyCQYjHOBRWrpgFhVDZUcx9IppQBiwt/0
mazw/zxnFNnLQEyDUrZlK7lAoFZf2fVESEgnZiOD0e2Wb6sN9vJriC8EJch7ugvi
QnVfVPIfyNeOdQVSZ3ji7LpCKRM9kWohsXYGMNIae8lVvFU+a1pfmW6Bg+PQd4PM
1ECReLeiAZ6pu5+fQgkEcfdAkGpozUijGsx0kv1ZdV6n+500O3XR4ZWIBjNf6q7K
CH/I2ck04CGt0K1TtRhhz4E8NDbXBVtNYLztBnFx4+CH84K7C9JkhN79m83h8U8b
CNHOtKdRNFO/mfPZCilSL8Nb39wLDol7L7zOykmYIbI=
`pragma protect end_protected
