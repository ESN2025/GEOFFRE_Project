��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:�1A��"i�	�x U��p	iԍ�Nv�l��˥A��Hr��4v\��9�Pq��K�6-�Ip��s��D0	�<�x2�"lŔ�Z�� ���#����{vEu��ӢO��#�I��P�!��'����N��؁���/=�4>hCN#����}�P[�O�Cޏa~����F�9��}&)��Ʉ����{�G.)���˩�ql7DՎ�S�N�Gj`�ge�H����z�󤄺��E~�{�`"b�	�^)rW���(=��'.��G�wT���t�cDvcp&�_�gvF��{%%#z�҂�[��n��z�4�h�
ș��M�M��'*p���LM��ۤb�\�0�z�W8���N�v��<�f,��	ކV+�y`�A'�x��W��j�vu1.1�t��?Je�GmR���r$�/)V����QeC�e��"�zO�s1Qq�M��y�,�����0
�n����,�Ir0SK7��9H#�E���+k0����3����@��ȗ�"5Y��uRS���!�_�!�{ø_��B���L���K��e�T�����3�����9W�-�����v�T��Pm����|� $-I`���u�bq�����M}Jj ӗ �|$i�Y{�#S{@N
Yݹ6ʹ$���Q�5�3M%\M�/�<G�oI�,�Q(��Iu��~�%�(�����g���9A�Prcݜ,2a!�T��L��	5A"�87w[�t�kP=ԺK\|�d���3����n���[��g���!��>tX?� �������	P$�#��71��9fu�p���h˳[[��f~I�I���Cf��~u_]Z�E2eNd�G�uJ��gH]���4��� ?�܎�6����m�8��3�	����fkr���阚�	�P����u�'r9s߅{c��nWv�;|��f���K���V���Mq;����u0���%=TQ��p	�qwߓ�J�ծ�a��[���"R�Ё��T[�e�t��6�"M,Ȕ�g"ǜ�\��&��T��J���b�$4��f�b��é's]�çCH�U�oޮ�G� kc����Չ�s�������؄�����MP�$. ��2Kv���kt�_T2�E�]ՠ�s��dQ�������@ݻX��W��"wʕ %�;4H��S��*�����^��^���
J��iU-H�1$,Z�G��p�V��۠�`�����YΪ����DvK2��W��c�����o8ݯ^�Tvw3�(R��tW�����/�#_h�*c����+x@���8aCG�Fx�a��l�Xy�9_���!=�x*���;�D���_�dW��E +vJ)<,�feF�WY��[�lV���d�1������k���v\��?�@�6�W�yg4jl����;��A�ao��.�{`Wc�����w�F"���,5v��M"t�j�+F���c���}�a��}�z*�þ	�+}ۺ��V��0({k��4�w��D�4���1��T�?��jQ�Sk���bU�_����:��Y���9\��Os�XV�KWn�}�RA��P,���i��]������J�T/h�G�苖���<Yl���i��`G�
{^�\�]�yje����A�:|�;�G8K/����w#B<� J�1H%�p��
c��^�Dڕ�\���4e~�-�]����A�B�4��o�Vj��kL�R��$��@��%I�g�?�ݻ�D[pҌ0;��~RJ>'������Y�E�'4Vp�VF�$.�+��6������'����h��%\p�%�̂����0]�9�|n�$w����[���ߜ����Mk� <JP�#G�nT���7�غ.~��򷶁�s��|c[;v�_�[޻���n�.#���h�4�5��(Cb&�r(YW�nM�ۂ��+C���Q<ߞKY��e�Q�<�Tp��ū2̧�SODLk�/��
l��7��N6_>g�T��IJ(IɅ�w2�Z��{?E9�B�b���eLm��I^W���rF�,��N��.ڑB�Z�{J��D��.!�z�:�������@-0s�l�v���~;/QYɸ�O�X|6�C��|�h�g	YT�ЅI��ѹ��A}�	�o���y��	�m�NDE���C�A��14���P\�<L���k�{eߕ�e�Ԓ?�2�R��an>ќ����eLC����%I�-�轡�W�G�^2Y��h d��"$5�#�&!S�ىa�s�%e��u�8b��|10RO�g)���p�LO��R�;�l�%�~+����b	3[W(?TKD������
��q�a�$�����:�_m�]p�7���)�E�]��*�e]��OJ�?@M_DVN��$�)&�^�_y2	���T1��'�_G��Bq���cj@A���m0'?p�]\wG�nqY[�nHlWL7ߏ�z�/��}�a'ѝ�Цt�
?��B�������4{����@�e7о/B�g��	p��jE�n#V�G��:�L$Z�؏2'��,HEǖ��p���6O�����l���bҝ�iG�)�\��u�i�X4���a�Mz+H��"� ��t�YC�`�%��tXüg:#���Kn��������
�$����\�r1�l�PKT�aӴJTP#�Aba�.��c"�<����8}e�����	9�r;6� �ˏ2���<�1�x�b��{\��w< :�ϢE|tGH�I��,�π�]/��<&0���a���S�$�c��}�5�-w*�z|Ȑ ��;�F���-���g����]֐w�N�	�_�������_]A�%�iUz�L.�A&j��B�q]%��h5)�����~φ�S�<��W.2�	�0����Ce[ �r�]i��V~J�,eP5�,!CX5���h�Ǳ�Z�Jx�?ٍ��u���ބ�F���%@����o���k#�0��HNj�'2�8���+ֵD%�6�=��iC��"�ƞe�=�oQS��+o#O���	������''��y�jrY���O>�v
���M����J�r񳉧9>����j3y�#�Hׇ7f�u�d�&Z��p�Z���J�ǧ,G��h\��y��)����i.ehjZ��k��
�&�h�ŭG�</j�%�~�� ff8��*�<~av��gh(��"!�D��`S���xML�1�V��\'sH_]x��b�˂�䠱y��w�֗���ce��G!q�Ex���t�k�6��Ϣ Q-r�UD~.2N&�5��ݬ���.�>�)�?�VGh.�^  ,)����j�z^���o�sRQ��ߌ��aQ� �X�Jx��e� %�� #)��/!~�P."���+�;p��*r�TY��d�eVSV��ƌ���É:�l�E��1,@�Ȳ�mC�H�&�M*��S�>�\�gd?� Q���6NQ����k�>{�����6 ���R�XیoǌLu�i¹_��l�C�x�-���oR�C ��
�"��/��V�h���윽��X,�|�".%��u#'F�o�@��mJ��&�q�vR�w)��xP���.r'�����p���s��g��=�z_��=�����<��$hv/N>s���d��2�N��ח�[O�ԓY�s��[��U�7n 7`���U(���+D_���"�s��t���^�K��P�)DT9:����Fd��'�(��+T�S|
Fg�ig���E�P���B����P�w��|� "�#C���߫YBU�j]x�94o�M.aV̼�-0�wF�	`A�-�X����%d�ݗ�ⳅ����f�����ѥ��y��UO��CC�,��ty�]Ƒ��8"T/z�DQx�����t����'8��0$+���O��T�К|�y��6��FU��#x0<���2�`<���/��u,�oY#���%HKF�jFROs���@�i��Z�LD��J���{�`Ά?J�������s�͕��?n'��4ж>c���R���u�[��(0�m��5���� B[�*��h��sj�P,��	���`K�j�[xy�u���|,������~�F�|��U�����'G�`G���^�^��f�5~��պ�[�Ey�x(^C���e�y����ATbq�%��V�mS_u�'t�}#�����>�\�+k��"�I){�4���㌝>��
i�/����V�f�u��!�6^��Z���B�����˝�v/)&� �i���cb�{�5�w�
�]́'�k ~Z��Z���	ls��|�GagZ��>��Ai-�M�@�\�x\��$J �L�rh�9O������K�8�a�~��2}����A����@.ز�����`�:I����5>�}(��|4Sw5�S�ʔ�������i�����5V��)��Q�-�0:��)�X��Y5h�d%XZ��������s�ܣ��okO>��fݶ����1ZuA��s4��1�{rXݾ��.52���V2A��$�!%w')����@�yu�?h\�lWlʕG��7ʑ<�'d�d7��|O�\1�׊޴�1�c��b���.+��F����O���F�%-��֖��s4Nb��^�o(�X~b��������$���>�=�R�<�Xr{?§GÐ{
�7�D6ک5��@V�D���ܖj����l6f��L�Z��"su)�ͥ|G5�Uߑ�W�hX%�Q#A��_x0T�t7}k�����`;��	��Gd;elCo��67��m��@����H�mg�
6�ȓ��F��+�M^�\[db��}b|͏f8a��/c�V�K�C0�ͅӐ�Ǳ>�+������'p�34�cZ�s��^�y�ګ}i��fL��`T�����k�:XO@���NeS_��C����!����Q@��ًb���Xu_���Bk2�v� Q�L��[��n�z1Q� '00F��I�q�d�(
�����$fO�����E�)vEo����u3L��l�>:5�A<����|v��/��3�g��E9H���L�]i+��zu�s7D--����rOoY��!.(�?��ƙ�)�X�P�\�7�%м�v�ƮĠ10���F�~E5g�*��Z?���� �/p��({���;�:����`-�
�b����/�F��k��,��א0D��ɵ�j��23�a�ŵ�N��@r�=�o+�¬Ď�`�];�h�po�m��*$�k�")����^� N$�\�:��;5��kn�����0�a�d���]���Fg�w&Y�{�[�uڭr!&�hE[,!nۓ^���,��X"�Qe�Փ|��޷V%�_�Q8�=9-�ny~싥H�ѕY��v�52�Dbe���_h���J�Q��u�#��[����ָ�iaf�cR��>Hm�_�̸�t�2z�L�^��`{�4�8�Ja�Z�?���o���ZX)��Ps5A��J����J�������ѳ^��"��
[x�)|.�D40-O�d��j}�$�B�8����ɥ>�׼�ʌ?{_'_[�_G���	�+@������u��2 Y��-(�uu1��W�4��L�Si�$��2ײ}m :�w��h>�`_H����b�}��3(��4�1Ng2V�L��q�kM�t Ff���<26�!t��fgC�=�:$�&�5���O��A!n�������|���aq׽�0��c��Jj�θ��q������M9!���t��&#9��@w��W$ʑ|�|�����x!w�C��Ç��>�n�]��`���Zr�!�JKн-隍��KD����%%����fO%b\rӡ�x��ŉ?Gi͞Y�.܈!����ѝ��8/����F�G��]��s�����w�� �[=a	KȍD9�ֺ�Ї\�`[��8����QJ�x��1�n�������(�}�6��5�8�ɒB��i� "�{�Q�v���J��gcЗ��UJ,�D���r�C���)�F?��5�iķV��')�
�?/�Uzv��^����Ɍ��Tp��,k��8ݓ'~�S9K,$pF�9�����t,���"��q����@�w~/DGhc�c$���q��.҃6����A#5{S}k��%�6����:$����[��"Wz%�F�����?�3��"��(�b��*E���"g��2'=���œ��ѹ�P<=�ukrS��������� ��g|.��Q�҄�f�u��'�U��3l|�YBv���؞�-Ґ����,�{cw�O�O <����;|��:>�	7��viM��G�F��� ��i����D�_�_cBψ�LL7�B-��o������B����Axr�.�x*^�:��B6��@s>+��Ө����c��ћ[�`1��ڥ���K�yXe!�{B�q���{�̫�Ȝ2�9a��'���u�ե����L�>(�8�~�i�'��R����]�u�4��K{�w�����X1�����s���`��ىl�'~nO��N�츮RK����n'����e,~q`���b�����E?�O�?��I���T�� !�2g�� Vb����0���9�ļ��5�&n������_G�i��BY��(�b�����q�͚���������R ���q`f�Xv� Oo��ey��eY���k'���j)<�(����41�$U:�	b;�,�N��D�'���z�2ꗦ� ���U�se��Ef��@~6�P��#'�&l��;�դ��.�C��x�ج�{�����yg�o|�vkf�`U�ls�1��0�VĘH�5�|!��dA��#T��c��D�ߎ��X�vyXڨ�AW�c�O-�b�idȷs�ء;���V<~b8��x�P���c�Z�y5�>�1��0�j�� fl__\c�2i�tmC
M)�g!-���^l���-eT�e�p�GA���3Px �~�������w>��#�k[¾�\oh��z9�m�H� ��^ϒ5X�	-GU��
7VMPL(%��z��a�9��a�����k�am����"p��q��y6'1>�l��%�ҍ�,b�\����۸�eo�#L�-�"RBq�����g�M����M}}$��L�ۥS�-�y��4�e(dレ^�1�.Ӣ0Ɨ��x�dN�P1�R��,V�S�z�c�n~�}�8���m ����L����U�s0�D�����UΏ���b��ӱ?Bhj`�xƮ��w�aܵ�U�b�Uz���c뢲�����D���6cN�t^I��,��N}`�rv�`�P���-����Ɩ9i�`]0F�q�Ϲ�����cW���[�)MO�P)�?զ�{����:m��k�&.�VOe;G������!K� ��3O"z�@<yBVZF�f��5c;�g��ACB�����}�|$���K҅�4$&���k����zXS��R�T�h�#�U2vC���Wꖒ�w\��U���<�U�Wl�G�Z/#�ofX:�gDS�[�t�	p����{:�����%�1��7��W-�c�H��H�t�aVBD��L������z)�n��T�U�3D����I
c��n{�bb&���\���4��PW�`TD�KY��%.���:p	^�Z�x1;�ݏ�����{*u��8�*ܚ21<�Hҟ�;����er��T�����A��O"k`c�f�W,ر��c��"4M�ou�.�4�V�pVϷl�fu��a����fvr�Q��=�4�pw�En�~,��j'S�.���	a�H�	H�a�v)���F���q~����f���+D���??H
��Ga*��p$l��D[��p)[��=�8P,�OR@�b��1ܣ���jg�d�O�r&�9��#N��":a�`�s�'��>*�Bf���*m���j�d�Ƣ��^B�&W���[w2�";>#ENw��ꊶHu��v�/�`׍h�lz3N_�c� �^��=̆M����@�l[Ê��b�-쾦w�&Ȍ�W]��d����k �Gc4�ew����i:���@"�ne�d�i<wY�ٗ��j�:�o����~SX�$|FI��D��Q�/�oJ���;,�M ��:�z����*��R���$�������2�{풌�0د���EB��6���LD��H��iD;�0C\�?{W��$�ɦ�s/#���8׷�L
9�.:бi������cO���گ��D�l�2�gJ���M��*��`=��O�'�����  F d́��.ӕ " �N;����A=�"���������CpA_��4���e��q0�f�<k�a�74�n~P+�3n�|�?N��瀔ۯa��ƅ#��4��DD���pc#c<�z�W�v�^�En�yg��6%��x}��҂��J�'_�J���i���J?�̌��=ɾ����+d��GR`Y�숋'߽��/�.2��eB0Ʒ���������áa�oG�Sģ.���z	k���b�t{ݠ��{��Pw*��D���.ۧz��h&�킑#���'2W�L�g8��[���Aq.5wT-�)L�"����������͑�j-��3��b�I]����xk��(�������HU0s���߲SOK
� �i
2`2�$����B�+|���>�:2:�N�*���1����]ov)�5 ;3/��W��=��l�VҼ#&1�|��e�;D���Ň���n�l?�YI��?��g�����2>�?� ��N�#^��]�B3H���8�sI·�Q)�z������U�>Xم�����-޽q{���+��1M��/�\�E��X�<�3\��Y�:�/O׈q�}o~�ZGۋ���ij~��oōB���c����l�O�e?��蔇X�L>��xB#��=��������?4�~G��]���3�O�l?�	�I1~������J0W���C_d��`ݯ����̲O��^�a��Sv�$���B$_��ʣs{=wH������d }E�bC��MN��̜&e�Hxz쒎��	��1�|�.U�W��_\2�����Z��;-�����NO�O���j�{�ݸ�PZ^�۴G�a\���X�j�NL�g�ٛ���yT@1r�5��$ty࿊��t�f�8�j�3��)�w2)�>����=�K����wѰ9�,���h�%�?7��U�!Dr�5
4�P��T�����n7$	��ۉ��d|G�oy�-z���0��&F*Ȇ.���,��`ȱ�t�i�Q�0�kV��|^�P��4KR�E����,?�³�^҉���'����=D�(s#�$��	k�>�a1��?�؊5��h`4[{�V2LǷ]�U��S136��Q��B�.>�-�ZD@"�LY[�`J|:��N�?�My/L3��c�E�G,5���<��ln��h��,��e��.��[��$�2Ky�7��Y�J��<��Q�.���m0C�9�JI�G4#v�YVAɿQ�fc��]7W��b?Wr8t<��&��A��L���Z.5Kb��Ḱ��\�lXT��l"�����ݐ�v�e'�>�A���hX�9f�p��k�!� R㬑k�g;wmQ �5%�ܼ4����Ǵ�yh��"	A���Ս*��.��U��d��h�Mu����y�i�j��1#}UeY���+$��k�^���_�,xB&y�UΖ_���&�"'�$�M��h����7eo#&}���A��a2���A/U��h�h�j�R�/����v���?��T���~��ȡ��;���xSqo�)6*C�vh�J�\�GK
r� 7 ��!���]Xe�%o�N�'�ӓˑ��5@�[U�FNz�
��ֿ�?(���]��/oHc!�������P��M�]�s&��y��������Ҷg��j'6t�&��Q}���[+���b��c�c��K5����>�Ua��<��E�Y�;@��FEcL'��Ѻ�w"�G�{��_6$7&h���!��8�4�#F������'�|T�A�o���ghuN�t7�R���ƿ.���6�=/��|��ºH�������W�5� H�1��N`�(&r�5�粗����ԗ��g�<�w�����bX��9soz�\UG��	]Z��҈����Fc�}Kf��>[����k-�F�h�~��%��T�HY��UJ�I��%�/��c�� ?4K�;��Xճ��]I)V6�t�q1� Jk��W��H��*�k|��d�r�3H�ӣ�F���dm�T�>ܽ�o�e|�d~��/]��sdL��=�]���E����.��Wc��9+
E(�7�th����"����=��z��J@���Kw��a�C�K\��5�C���*��ӺV���68�5�t�R5;O'��,5tXvky,m}8f�)�m�
O�OƬ}lR���2+��T�$o-0'��^-�}p�4idx?cT��e��O̍M	�+Uy�x��R��'�!�-ϻ��a>�
�0�@�@aQlyG>�}ȭ6�|�`l��1O��r~!S�"�G��SJ���2̙�����U~�}e�x�H���oo�h�2ê>=��1������f8%�͝�f4�2|�2p/��|����a��W�������D���d�q�ë:"W�x���n%O �u�c��1�*�B����7��a����}�iѻ"ְ(Z�K�̍�_�ce(�_/�񖒞��Q��ӹ��&z9C�{[~�#+�$_�զԣ��2�#�F��� �X�V�f�,+�om3����t!:�&a�'����_���C�J� 4��B�;j�ʬ�D{Nd3�{�]1�W�L����i�;�RFt���t	�I��.�����3�H�@�kX�E_��\zG�"ED&��O��$���2<��Kc$��M_�{.����	]���P�o؛�oꗶϳ�[,q֨2��LL�Fж�Mm֣��aqN�s	/�������"9���^��dͿ�9Ǔ��pL�Bcݳ�4�gǮ]�"2��/W�/�h�BX�}�(Ք����u�wQ�
��k鼃^h��X[Z8.4��ӆd�C�9���ڼ��|�8<�1�Z%F�e$�Ϣs����z�T�М�p��I�X&Q������� ]x��pE���qky}[��.	��j ���w��w0.durS�X���%%V�S�ǅ�P8P��T�-�����]����kA�5�q�e4�j认�������`�F���4f6L�c"�Ǖ#Y�{=�)��[e�e�����W)LB���kt_}"�$$R3߿��		�O����L��pZS�}��y6�n� O{���|4�
�@:���H���g�RU��^Vu�����|�@�<YZQ��q�c�YuH'�x�sb [sd�%8<t�Ae<�<������M��B/�+� (��E�.��!�}��Bܿha.����[����C����t�9HQ]9�}�M��O��Gsz���w6D������t��Bj��� �Xi4 q�2c#+��1�Z:oK�f-�r�p�Al���i��.Ė �*ە-��5���l�q�iL����b��!���^V�,�>>�*��mT�Z��,��uL��w�U�(����	r��.��xS�&,����<Å@���q졘1�i��'��?�@䭟ˍZ�*����;�0�}�
*F7ᴈ-5��l��՛õ7�!�d;S; 7�� ��j8DO���*���ŵ`���^��;;(#8�Obp�6�]]����sS�A�8�������j%x��/1=zq�cp|R��;&f,��>=톋Ff*���e��Ȭ8�9ɷ�J����-�6�Yi��q/*��`@9�=.�i��p/���"�Ȋv܋���Yd��3�0Wd�Ζʠ�Q1�o�,����\�����N��A���?֛~&����\�A0�O��b�O(���}����'e�1&
��uU���3fs,��lN���`����H7��izԆ�K�wtDF�ģ���%߉�l�cYv򝩗��F�`�}� F��4M�r^��bht���׏FA�Кc��L�	�������x�՚̘�I߾��ju���N�j�{�5*�1�}�B�$�}��h0�\?t�*��݀����{.�ڢ�Ak�_���(S����(0$�	TBZ��K@th�VZ9O/���'KD@�f
�kϡ�3Kٰ��l&Z������R��SSv8�{��:��
T��
�0Ȱ��R�I�ۮ��	�W}��ڔUy�mf������f21�v�
��o���9�"��Yg�i��7a�P�V������ߍL�����нHb��<�秋�|M���qC��u����;	�B�wΙ^Y���g_����~���z򙚹@��HDâ����-y�J\����1:����@�x���ҎC���ciy�������-D��O ���"��&�x�|	3p��~��rf	e�?=NE�E��u�!Ȯ�J��N8$_	�St�@�iѦ��BlX"H��fY���G��=��x���B�j�S��� n�(�?F�+���)⫂��0ێ��G'�qdЇ�0N_��6�>l���s,�3�$,����ز�&0VD^����@�z�*�Y:���(�_�[�(�n��N��ƙ�iGT���R_�F:	IQt	7��*�E�za���-�J�������P�O���6dGt�ŉ���N&��%�J.��%˨zI�������Q�2Z�e�2�F��W�c6��Mp�j�-��K�/��Å��i��-!�K�m�L;��:i��;=8䑗���@6x��2pN8�<��B���_1l�����$�c���%k����5��T[_�0��5���K�RH�����a,���(ѹ�}�[��&�嫄}c�31�ʤj"=&��c�_��OdW�.=;�=���"���F}��H%o��h����9�U�;�X�
�f�+Rr5i�0�^�n[oA���sM%';���!*��6�X��*m�Eq����9�Ќx��,�|Vl����1 ��4��#!Y8��'=���9�U��ɯ��\̒��{��%
:���������uW}V�����-�N1oˢ�w��.�}
U��nR���I�~ ���Q���`���a��=��8B]ix��������pg�1����P*�M���A>$҉A�~x�y��3��4���Ybݖ�	���O���@��e�uΛ��Z��8 �g��#�&GS�l��}Y��]h��"iҾ���5W�-Ow3�G����kH>7X�>�-�������g�^�RK����� 	�1t�|8�z���Hˢ)����N�x<��N��q�F��+F���/������Ո�I���@pm�k6y*�N6�fo6l	���c�bp��]�k�I�,}�t]9�ò	[�A���y��׀5t�!�l?p��r5���♣;S2���a-�������-��JB��
w#3��E��p^h�ؒ�˼�`&�� ��پE(���[U�.��|'p�9�g���ܥ��i��0�6=���=��+�����J��[m�KϮn���(�k���s5�N=ad�Ǽ�	�+������Ą9��	.�bq'ż>��
���#��n+�R�4�1�j��mQ�*GU�c��]�Vȵ����r)%ܣ��[���m�U0p\:�#��R�7�iА*i�*�Vk��1�(a�Z�S��r���Jk�����5���s[m?6`º���u��n���}�5e�8!#Ur^Q�٣�ǫz_8�ъ�?����������:���6�*�yz�O~�]���	�1��0�5��Q�>Q���|���P����-Kn�z�plp*a^�8�~Hо�{�Ř��`���M�e�� ���j�ȵ�Ƕ7��by���#*.>��VIk*1٬����Zq G��_�c�Kt���O������%x08N�@���'�\�X�H�鱋���@�^ɀ�z��~r9��A��A�W�|u<�,2o��E��ݫojm�yb�g��U@����+��[�<��'����,:�Q���*�Uehe���-�cg��>eƐ7U՟B?j}�;�]q�
]'6�T���<P-�����ғP�g����#\�{�L@9�b�28��M���`��g̔��~� R���|݁ ^�\��O���MJ,����$�\}u4����<C��ݧʏuvYnk�9G>
���
������h���0��%3�k�h�'�٢�b#�Am��I��R[���eM7S/��JL��3}���.�P�&���䉱��'�v˘ۿe�R��_��S��7�]� P_�T�F��#B��_љ��S&(A/���O�k<�ҟ3�d�6����e�
۠BX&�|���ɺ�W�`��iA�2���R��h�:e@�g����QQ����U|�.��KX1����l_j����s=���Qr*�j.���~�5w���m�2�2�]�`�7`�@�0�o-���&C	UX�#�`O��F+3��m���,���3�Y%tݲ>�0�P]�5gȤ��
�y�!���gWż�P�&�:h���\jf�@5Δ�J߈�M��Q� q�܆��A9 ���gP���iT��H)ʰ�~_x	�۪a��]��1k���n�1ĩ�����5]�λ.o�GL�)\�e�a�@Z�u_ �~�o����l�Ń���Zf�*<=�w����hm
>��Y�8�`{Z+��"_8"��×�iӨ��rB��!@�}�uV��V��ﮣ�N�-l.��� �(�n�2�ʰ����:Ô��OL�W���#jT�+�����
e��2*����W���/T�{6cp�3�Gj��YD9� �hZ�<8=��W��LV,yC�З��'.���p o�|ST�%:8%����o��+�̕���i�V����P�qʺK���s$�!����e����v�	[Vi�).9�[��GӋ�{�֯x�}�Q���L�n�3���]�f
v���K�Y�ȉ�ײ̆�����H(����x1�����쵨�Da5l�a�V�%^�@�6BqV< 4M�������C܁w�]�qot(��`(mLX�JW����>����y���6�^�p��%�|`���k���@��;~cmJ}2%���~��7�+9�:D����$D	uz>1Ͼ�kܵ@�o��g%F�'t&��r�!�G���R�7�n���fɿu��*;:�d=�Ǜ�iEi���h��XMG~ n
�����z�v�e�y��-v��?���T���`7�4M>{-Xr��CT2@�0g �8�_�U�ae�!��Q����ǃHc�2@&ƙ\+lo�|y&�3�� ���/K�X��u7��3���3*Kg.yvR��\�p;���8�/�!*���-Gakyۭ
��(F�¬��M{�4Z���-į����,E�l{��az.G?iS����|s���II��M!���IJ�<`Z��<g�>j`	�8�$���p��ry_6����O��䑜0�v�=�< �=�l���?jbiLن�����Rx	T������o�z�j�Fj���=���,zb8����ma�j�sO��P�$j��G��7��h��1�v����_@�*}��t@'���# ^�`;���=�q	��D��l�; J���܁Iz�O��<=`�oݣ���
I[�A{lhA:=�a�GK��F*j�Fբ��M7CC1u����R���\)T�i1E�2��1r�^99�S��{ף�ݖ�D~@��d����HѹD .�m4'�m3a���~�A�e�A�EB�6��Π���Ov�a�tL#K�/��5z����Ҭ�8}@���(I��d�C,u�;����zW`ŏ��-Ԇ]KM��*v��e
.D \��K�hf��tN���ob�x�P��(jBY�X��Bٷ$3+��̚oQn)�㶹���kW%Ty��ʕB�m.�(ʹ����ȷ�$S�����	�����w�G�"�T3�aw��Q �v�άc#ڞrN��cM h`�_��n���q�� Ň�)?�`�mW�x4��#�.�yQUId�}�I�o�L�Ja���p�_��	��[ ����,'�R0	��q�����~+�;W��{jz͜`�4&��\a�sLWA�OT̢��F��̪�j<�(Ա�������~穑�w\M^C�2q��P҃!��5
�� ĳ|"x�VE��њ�O�=�w��t���{y]4��p��4�?z�k[���#��%�rr=��ғ��h���m���z4%9��!��H@�e��i�cc�=��J��7Z�����%X�W,q���]���gGhXЋx��8���ϐ>L�Bb0��h���O�Aa�;\��&��*�[��:�yPp����ԭ�ꔶDJ�6߀q�{xa��>��� O�틪����N(q����h��s|��n��T�1���f�H��bjt���␿	M���KhMu^�<!~����j�Fx0�:.��W�s��>�D�c��YҸ�O:#Ad�y<	DF&�°С'��PmU&E=���i���Wkh�3��3I+M�tkC}W'��Z��Bԫ�s*�"��\���M�[��`bѭ�
0�'͖I���<j�2 ����	����;9���
�7-�*.pV ~nz��/k�rI�h�։ز���y�jtj��&��g��+�7�A@��u�պ<���r���ϔ��v���S��K������e�9�،?���#�����g�G'& �q�1����'u����=U�<5)r+Mh�h��0 ?ӑH��>�,%é�TR���'Y�U����H�k���$_O�M���e:�|Ii���E~��(���{��w|���*/|����h��}�)mm��DIv��g�qe�M/�J����s�iF*��&[�$�N��[0�v`M���u<H�������/�ǿ���63L�ȇh`����=��Q�Lu���#����k<��a_TdC�x��$&�uLtR�(b��D �g���i߭D$��#�������JD�]���ٺ�xZDÁ�M/��e�i�t�E*8D�21˚� JY}��Mh�KgmhB�Aj�����	YL��`�q��Oz�B˩�e�����wfj=5	�P�
��ݘ��oRD~�%��\n�v����KLu�d����vF�E�f����m*Cq�%�r2|V�ԏt�AU�Ahp�w�#v$oc87s���98�:pf]G"8W.���Wp�g֑�Vo\F
E�67Wま9 ��(�j
`(������7��y��%�c����CP��o�Z�P��aDI�l
:?/k���H�հA<ŭ�A������1��&�%�����nTx{��6���|�?iW%�R*.1���(��@k1,�����}��Z�`5d�M��Y�BD)��2S�4���g�V�2ԗ�8<D
6Y	r��ȂMJ���:�9����L�1 �����,�s$�*$�t�6��>etX�DS2�n��ཆ�oJ6�	8z�`j	#�C1�/�	\�%Ґ����}��1�T���z����u�X0�Ձ�R"{n#Ly7�5���fA��Rlc�r����8�����
���`p�ƖRƽp�^���ή����RƳKx��p�� :��Ψ�8�76���A>����� h��O㬌̋����o�:��c��/K�yq��m�I�S��[��1���:s��o:��5V��b��&�	�	'}^?���;v��l�؎�)�j�6f�r�C����~���(Z>T��$LP؉�0�_X���}�3�fHȃσ�NF#k����X#^������@��ƫ�_U�$���;L��GC��s�_���7�7�KCN���_��C\p�Y�+��M��_tFX��=Px�nA�����5|���H[�Gz���ħqO���Аz�'��'Pדb�<d��� DVN��<�V&r�j�������tja�l��w�Ti�n��$�R>�@��-�Ƥp�=&��H������i_k�ұ��c���3��?���9�1���#�NTgpE走�� ��U�4D�e"/c�jdt�)��,�d�H��טt"�	�]��3R5W��GNа�+����g˃�{�y�Q:r/_U���{R]�Plۨ�K1-���(�=�A����L���iE(�G�Us3�L�Ʉ5�,~V��,*c��2|������wP��W��ߘ����Į��d�r�}��\����o�T���k�.��P���+)*6�D4J��0F��@|']x���f�kO��'���K��쏄����<@�s�C�3�fɲ��g���ίJD��"�㮣�Q����/�(���s]�R)wI ���ǻ�S���>[�O��L1Ë5��*q]���m��`VQ3�^7�\��E1ў�j�?��𭾑μy��<Tlλ8��!(Tl���%�k���"�Ч#�Kf�p'/����~�&�[u��v��PQ-�[)T�� �m�N���l�F�\��T�f�B�fu��Z���u�+Z�Cl�k
� 7ОZ��JPuC��A��?���w��*�To��H�1���O�t�I�����r��ؼ��+"���i	�tر���:���2����p햼��F
 ��W��n	�0�6ylð��{![�
��4e$�_=9pU\��McFߟ�w�j�A�Xe�����J�ܓ@t�E�� c������&��ŠY��XT�'����B���o�"U��:��q����b��2Z�hp�$����U��((.8M�����������|�Xq�ݷ�k���'�Q=�P�i��&�<��5G��Zyܝ��O�2�/\�3����"L��'fp�T4>�_�j�zL��H%؋R�k��(_��7lJH�K��vI�o�.�d�-�%���c܉������ئ:��ދj}�3������$�c�:�E�N{PR�J����Ǖ4��j������oRr�8)ֲ�����M��R,�����3�᎓8>Q���S��F���6�i�]��[*��w�J<9��꣯�b4���� �8b m�U�oy��:*��z)h���[ۢ����]� ��`�K�����D/>
	��"pH�:���	�kW0����g��O����7�?u����KT��[�s!���X��}G.q�2Ր�����Vi��r4%O$�����ș+]�{0�)��ۀx}k��}c�?,�<~�!�o�[MRyg��̒�k��UWΠ�j�)�q��t��P������|��w<O�귅��,�;A��9��ۨ��c��ohVZʾ7�I��]�r+��&�Rm��$zٚ�o�Z���K�7�b�C�ɳV���/]c�0��:O��H��uH�i	jN&��G=�홹PjH[��\�AMs+xd�Mq�E�{5.2�B{��ygdҖF�1�T�=�r��w g�N�ҕt�Y��&��r�� @bce'4�E�����jK{,��_�˚�^�-U/.B��L����__,|��yuT>��h��('��1����x��Rϻk��PLf���Pg�]5NВ�^L(���rD�I\1�ܞg?[_5�ZV�G�YǯH�&���4�ug9bq��Rvdޅ ���0U����y��5�C��G���k��\µ�ʈ��;�X9i��߰��Q|ug�=�Wx�M3���s�r$����oI%�a��} �:����d�Q
Ͱnn?��vS��w*{����+���}㲏o��P>%����L�d�%�#���u����똩Ͽ�	����gy�}Ź���i����s������� �'	��Ļ���1x���*S6��+Ĩmf]ǥ���^vVlv&'�C�}�{t�^oExb �%0L>�4�$)`:H�$�*�.\Y���>K��>��<�;�c�b�c���D�˳^� ��a���C�`�.�
�80�� |sE��6\�T�����b�P���?&��/�ٱ���w���U�r�9�Zħ4�/�0�����b#�}V�ѐ��t�I7�T�t4�Y�}�Qs�6�	�l���D�T��c��t�aK~-�K����y�Q1���2i����N�z����������z$Q���j�@/i	95?3^��]2{������uk�wz�R��k��'�����X}c�J�3�ѹ�A�Q���zz�º"�;�L������iz�O�m�g�?
}�h���1� +F�
�����Z��`.��%�Q�!\�GJp��B�Z�Bըu��u�4����'ݐ,�v��2w%l@޽������f�4l�M#H�*;TD�P��.O����-	�i���}[����rh�LJ��/��$�2�'P陪lϹ�{�&�t�#�P��R�pS"����\�]�?���t;k����H�P2$�����x*���Y�{�y�X?���=;8�Yd�Ï%u�ٙ,�@�sA�����EVK�l�tX\( ��\1��ej��99ZØ1+�O���V�(������i�h��NN��� �f0Gg�=�oWY���xL�H�l���-���nMX�:MD�ȍ�Q�2bc�<�X�~�tid�4��jۭ�%.MH�*ء�� �!]�A�*���L
"H}��u��B(˴8����kZb�ҏ�7��M�3��ֵ$gW��a�:���ҡة�c �V徛j�r���,X���O��^}�Z��lЖA������*\�p��&�4/�;ε��٥���u�+��L�A9}�R�����TC?[+�^H=e�?�_Ҋ�^:�T��6��Hxt/��)��y�����`c�=��@rt��8�(�X�lƌ#�r��(�4�n��#�*�i�ƪ���Jٓ6�8e��5��ى�dN�r�#�] !�q��j�����w*l��~�H��Օ�%Ű<fIU+j�Zv׌�{�t��jQU��f�({O �O�P��������;�hO�8�4��}n��/ނ��w���ɼH��b�{=�n��ã~r����數����~��\�X�[9l�C_bE�j�c�P� �n� x\pFD�598;�|�[W���G�H�=��FF��"���j�q\ ��[Aɮo�1���Nnu6�c�_��{: � k����2Go+��Dr;��]���4�� m�НF�Ζ����֌܆W{<m����/@����rH%T�\��$�9]����R��tL(+�d���NV	lGr��S�=�#�Q�!c$��V��2�K�p��F���>b#)�����SVl���,d��w�k�R�5}{��P<9�;�߮ueS��	!�<i��mB�j��)��bu�f�]q��z�v�b7}�
��+�$�ż.T �L�qߙ�~}�C_�?�*65znv�C�2)��aC�??��1=D�d�׉��p��Ȣ�{o�B���1ԕ]r1j�c{���]�O�.x��@�J!A����;�k!/9���+�+�¶��+�dт���^�2T�����*:�3RU��i�n������K|����u�8�o�=�Z:hr�YE8@6���5�������v� 
����w�/._�]^��r����P�ٞ�&3�$�AQ�j���tsl�#���Q*�uQ��Mr�H@�AsE9���P,ldS�-7�x��� �v��������L�(��溝
�8�O���x)��xm���FK[�^��x>LٯY��ۯ{��I��]�Ow�������T���*�o{/���B�W�pw!p�R>��u��;�5��� ɳ5,���~�P������}�/+P���">w��i-�N~�q'ќ���b(�:���v�8�DW��Lt�%��4i�Q�)����$9�(��9���u�j���Aӭ�^n�&r�-]g����u�"��5Tf�<�I�&��]�P'�t}����O!�y�}���hԪZ#�8�:&�{�վEˢ{	�CT���m��/�˻����;�5Zl��kM�2Ȑ�Z���O^M�]�O��g�QK<�<����eݹ�ʜ��;��㊘7{�i�h0�z��g��vr@:ڛ��$��G���G(t��UqJ1�Q,�g8�&��������3�0�	I�������['xF� 3"�`�J��c����6f�Jb������P]V�e�gZ@B���&X��\��ҵ�:Vpm��j�9X�ǖ$(�М�Sg�eS�dw�;J��"�P� �!/��ٵ�\5W�/�A�3_��G�����椫!�c��2��B��F��p܁��u]�X�%����W�����5�~h�#V8Y�	1�ĸ��Re�Ča23��Z�a ;D������t4��<�
V�uh3��;��|��smځj�\��Y����,*c���+�h�dF�U��zlzZ��%{��<]M���n���-Q@-ރ7+�R���e���t\T�|M~i�����Lt�MI�����]�Չ��Szw���1p3̸��[����4���MNJ�mͪJ*A�V�{7�#��v	�[X����5�����yL7D����-��^~F�h������W�C��,q��Q�<��4TGE����Ks$Ͻ�����N�Թp�3^^�k�j�n�d����=2Z�I�\>���2��
���;
��c.�wY��p|�9q���&qC[lR�g9X�uw����|�#d{˿�{��d���!�8�ųk���S������hvWsH���"/��U��[AN��3�ְ��~�UyT������V9�H�2�h�D�]q������?�b��N�p~��(��uQ�ԜfmFߐ�����0H���֣�}�H�vz�)�&���x5�ҘC���q$��$��f��vg����A�w2xf䈬��m�\ĝID�/x\�����D��;t��Mw������j�g��I�G�&@9�3M;� 3��q����Zm�Yh�T+��Ρ_A���5_G�~oe��CnZ��K��1��z[3���q�W*ݞ,HA��n	���1a�u4g�Do�m�c/������~��љA������?�{`��m�̬=��wUG'c��u鞣�>�����T��Uͷn�L��U��d��~�W1��$�84�*������,m��;�bQ��.b����D�27���&���(7�YysOmF���jv<`N�v���Pii��]1��b�R��wf�&���c�Ȇ��_��F�^D���vC�����Q�z��+�jC�Q�;��"���[ܗ�p��;�Hk�	^o�4Ay,�X�s[f�����q�i�(r���Y�0X>���W�w`5��H2>��ԃ<�B�s�{f'@�|{׌��w+�29E/��Y��%3f,	)���*�r4�)�g'���@��,�����2��1�8���� ���~=:f�)_Kju�~�젋+��C.���SE�A��5���f'4�X /�u^݀�U׬G�ֈd�͔�Z��%� ">��n���ѫ[���I ���x�P��.G��h��xͶ�XƠ��z��A�F�d�7-�3�[���E�F?\�`��k9��p����J�s�(�� ��55��.��|p��+��]���<	0��	�3ȷ��+@z~k�ji|U����G��^����!�j�k���%@A�7����ޏB;��[�(C�-�Ҹ���˸��i�~�q��#��"Ȍ3s���c���W97VY����9�;�(�n
�Pȣ��8��x�s&�����j��;R��з�}#�Kx�b/,2��̆��z/�V5�&�#�"�5=Gt��b3 ʨ�\��_�]5�Zd�G0GEŦy_�Z��Eޣ����)H�[_�o�x�zSQľ�6ɧN���_��	+#��L5�]A�����q#.�
x.�ҭ�p�&������kP��Y��͸0�H����ԑ�tI�ؔV�-UC��I��n���:(��bx���g�\
tkZY������G�;�Dx֗$�:��-v!H��dg#v�t�)"��}����#_�9'5 �6��Ԓ��<�������6uu�~��cSJ������ZW���������J7��
r��E��J��Z��P/��X�Y��/��B����L��ńE[�
�%�����|��x~l5�\�Z=�.8rj���xu�θ6���w���A�xW��w�!�a��F_����8\<���q���$T%]��2�n�ʥ^j�/az��c�SJds��c�V�t�	_�4�Dke ���h����֖���%�E�&<��=�ǔ��Y�U��i_Ϩ?6�\ uJ���b1id��*f:\R�k�dg�����#�D���*,�z[5O�Pi�x���!5��k�F^��?.5<�Bo��~9Xӽ�9V�����g���O�w}XS}~�gE����zW��Y����=�	�><d�DFTK��t�-�Zfv��	�U��%0�!����r4������<�M�筬�٠�><@7�B�/X���v&e�E'�R�5�W:�W��4�n7��2�(C(p�5hk"	�y"��Ҫ6r�ja����\h�R�_ص_�����B�wQ����#P!u;Ңy�t�Zc���_���>�0�(q�s~-~���ړ_����.���m_�G ��]�#�F�"��o�Í�e����/�+�4"7�:�[����5��I��Ո��	�W
Po��m��ㅦ�+�|F|>��:���QO(��#�� �0�n꿒M�u�����H�haV@2��A}��zᥫ�!hE*8أݫ.	>'Ϡ��uT+Ϯ4M��X�Y��s�B��$UK?VZ2Q�^=J�w��կ{�9�2�E���\�@��X]f*
o9'�ؘw �.���
h���A�[8o[K��TZ3j{�'*��qP$2 .H榥��JA�ˊ�ז&6M��M(���Z���I,�ػ�����{�"p,��pRvR0m�_�`n6�I�v� +�����em^�Rv�p?`<3T���\N[zhL<����#w�m O9�M�[s�5G/AwƆ�v�N|�ǈ$��������#*�u_�����	$�3N�Vg��$�x�[�ô*^/ꇊe��%R_�݋���@L.�d�Z$�aԧnzo$�t��}
'�4r����KQ ��ɽ� o�	ٝF�֊Fu�pͿ�[IU7f~��{��"���3�ٔ��qZ��c��ۂH%�E�N#���-���R�'"�z
1wIN'���#�F�䜶�/�'�6�����I�-�[r{UGS�)G 'c���j��7����F�;�t�/l��x��:9����u��5t�@�	-�gs�G�BXʴ<��y}	���[��+N\��|�-�t�B����Ri�'5���j �>D�������]��&��5�/D��D�"Y$�9��y�#�z�+J�ּ̓�����qG�7�{��"Z�)\f��᚞�da|ӭKh��[T��n���Pa�����-���}X�cʑ�A����Ǒ�`�Q/ᨧPYp�����~�6�-	�tѧ����Y5��6�p��SJ!��*�d��<�Z���`��7>d&FR�g���O�����l\��
'�M�D9 �UJSd��f�~��%#�l��2ʋ�Hh%��]*�A��E�����$Y�8��u�'��MX�`�eև$�f~�-��0�n�iL���ia���,C��>�ûn:D,|^�q�ȔQ)������Rh9�����UO��L�g,*m�8?Zb���P`E1��_����
r%{'��X���x��w�2y�ݳ�Fq%�l��$;���?�� ӟ�F��e����+�Y
c?�Ճ7����<�Xago�����Ό<o�S��x_��W�yɈ��~J�o��6v�il�Rך�?�(yrIN��
�ފ���CL�&	3%Eˆ-�8��`�B����;a��PUٷ��}����B��QD��]��A/6�?���Cݭ�_��<&��s�>0wqi:�o��V���V���d2˙C���(-��z��d|r��~���1<߁!�(�������+��s�յd�`���B	���[�Us9�Av�yX���۱�g9��2��$��z1���gs�4��0cm��^h�ZB��Iڥ�o�C���c�����~4���Y���}�zS�`�Oe@_姍��Ζ��Ʌ�)���|SUe���^�M�k7�x���;� 9�f��ւ�Io�M�����~X�ڔkZN�'�� �y���شg�챱�Bu��,M����s�$�3t��)�n����{M9ӫ?l�G�����c$K�h<U�^�˯�.K���	E����uι?�Y���x��w��oX�χ����@ut=gR]L&��q�*:���z��o�5�SQ�5ʃ��{JJ�fZ��{�r��/v5
���:N�{؆��zJ׽�<�y#웺��̿܇�t�	!�!Q���T=���J��Rϧ�!y�72=��y��a��S�Y���fq~�?�U2R�}���sZ���n�-��+_�6`u�w��ݠw��s<��j�s��ʶr�5�b�W�J�#d�����A��ZX���v@�J�Qv��7w�7��t�:��+{o�/p�����\4�Vӥ�f�GQ�̷�,�Q�2�R��MBf b�(�p�ʶ����S� �l�:ʬ����ݦcGBE)�$���6Y�"����5*�����_�5+]OUG�B����q��^f��6�����:��U�$��E��P`QȄ0l�8�	�����v =[m(�_���|F�p�n��z������p��?n��_$[��F;�G����$֜F����ũ�,xqKg�L�}�NFexC�=�!�r�:��n���e1?N�'�)��D.|�'�)��M�}B5�I�j��:���D�lg��E�1f�p�����t�����*7���S4ga�-f;��
��D�:�"�3k].��
�X|��(�D���,�0P�n>�?�םk2��ٱ߷�=����R��4��3q����6�5���| y�n�F$fj��!�^��|}����<���fp\]�g^@����t�q���+T��q���;D.�1Eq8K�4�X�(�ҕ��5^�������(um��2h�
����nL��P ���ȱ�ǖ�(����K��MIL�����A:�`7�%%�� 6�^e���b(t��A(zK-(Z$���L��o���_������Xj�%��4z>�}��n�E�y�.0����
O&e���|p��.{o'Ж)�^�j�ne���}�d`R"���Q�yz?��l�����Jچb����+�]�#	saS������ ��V�r�D}�+���Zs��Ϯ�փ�C���D��9�G$��/!�p��0����&���M����טa����f%.�h�D-r�۷}�r	/d�!�7�)*�I3��6Ut?p�_p:6���� jO���p�ɩz����z;�QI�}[Qn���X�G`���ݛT+��0��&=��$���H��4�QF���,0XV��K�T�\=ύc$�����ʫ��ܼ���0s�j�}8T��Vߒʢn����e��$B�5�C�GM��'�`Pj	^�Sn����TѴ�L�,�8�SW����e�0����Z6�R����`fLy���-E"}�#���|_D�U!J΃�}���-sƝ�+m!�(D�O�1Us�<����D�@����ר�T-�����?�����<���_���l[����Օ&O .AR���C%�,�w?�W21}RzF �+~x� �f���h��}8�~R�w%��e����T�BOv�'Y���������%�@=����J���<��@JZe���y����l#�g�i�!�Z)�ƃ���z|��w�Z���& N[R�`a�>�<�/2�S@y��q�"N�� v/�
.h+�7'W�S��vq��V���� NV�i���C�wn�8��R�+̈�:��8��>���I��	gQw궥�ή��ώ�Ђ��\JU@�X��{����/�&"���a���.$N�9�_ڢ���O?�3+���"�ʿ�1��-%�e���+�1B��U����':na�f��� ���8���4���uV)5�xda:g~�OFBa�2͟cϷ)ۣP��������t���y����T��x�)�p|���	�iH�}b���w��w`��÷g��G(lC[�1�ǋ_i� ,�ە�A ��Swу�s����}t�s�j��-�P	+�M��YA����a�aV�]m�Dm��QM|"�(�[������m(���Q��M&"�@�!��'6ߴ��C�o���|݂ψW��Z���}M 7r��m_����EI��.8H�0X���μ|�uL��D�.e)i��N'��� �&m���|�F%����[d��}U�	#�M�
S2��qtG��o	@9�yG��Q޸��Ω����4k]���J����O$��������	�(d&AO=`L���k�yx����<*��(�6p\���o�� H���q��%澹Kk�*���j]7j��u��,��r�ve�E�X+���=FS{o7)uYl(�~��ٙ����B����O RO��i��ߔnb�ן���-�>�Ý%�Adr?!�ן�]sq��R�}J�竣y
��}�=�"��$�V�`ё�}E>7i���U,�XAV�# �Č٤͞N���e��k�wɛJS{u�x&6�!�K{6� 7�v`�3�/_��JtWQ�I��z� 6����"��V�g炐����N1|����@�����a|y�YP�&�<%�.74��8P4�����w��3B�ajd[;�MB�Շ̾~^�iO�#=�X����b� �-��{��:q�GG���,{�̄�/�I>3zZ�e����UO_ij.p|��zK��?4Y}JjU[F#y.�0A��F��j{���4Eo��4�І�"�d�MwZB�Mӯy� ��q!�7�6ʍԬ�L�w��"o/���4��3� �@�ղ��T��Qt�����VA�t���_2כK����O�!G��?ڒw��b�+w�(E�Y���=�������+�Tu�%1����t�ҁBt�fa~���?�M%|ki�M'FzC�F:*�;�0�K]��������E���k�0�`�]@R⯕�V����#ж���+?/2�P&w��"�^�,t�Z�:�G���ǫ�t���s��	�6K���*2
3��l����x>�P1z�M%�\s�)յ���]]�qN��ɟ���l���ܛ�؈���S��qWN;Q:-�Q.�6[݄!����<qZ���8�a�N���<Nl9��Rd��$w��#��+�z� 1:��r�D��8�.�\f�`�i`-=�[�1�U����R��o?�5"�2�f��z�W��&id��zx��@�[��7~"E+2��t���<N?/�=�p���E������=����#�%�ҁ����-�Ԅ��!7Y"�y} '�Q�Lx��S�:@��G�'3L�hM�_��*ꂜ��D~5z��^X�����k���]
֮�]�$}F�Z��:
n{)T���X2�dқ��
���������)�;�9I2�-`�b��2�<p+�]�� u C���{�5+-*�ƻ�
�RB�R�� 0)ִE��H���T�B�~�@�������.�2�x��� ���wM�O:bܞ�����x�?é��������$�X��F+�����p��Gٳ�N�i����bbّ=�I�������Y��|�?�.�;�X�40���p�|O�Q�ܕ�ݪ�Vs��~���T�̍.�7֨w�6̋������A������� �-�S8n�Ec��"D�C�z@	�JS��b�r	n���d!�4 г2�n���4�d�3��:ř97�j�K, ��~cw�c�����J�Xiv{����ٻ�@�8��bl���w�3��m�r�(�O�ٽ��]� �(<�4��b�;C��d�E��^Q����p�[��n �ԩ�A�R�����Y%j�R�	�;���N=Q���wl� ��I�+r�pR"��"��ϫÄ�pp�JTU�v�F��3$FŦ��f�I�C����a���o�x���U6����t���o5)X��C��~�y��n����[$X�+�V��?t�r�)g�z� �ti,��ڤE-=,����!4�K�O�U���(����ey���*L'�(�Sf�kʧ�l�7��_	S��z+Ӆ/v�(ZB���-�j��P �ײ�It�6�ՇH��"6��D��hG��3�k7�Tw)�+^$���/����x^��÷��=�-�O�1>A*@>/����z.�#�q������W\E';����=����%@�MUl���D��y�o/�^�J�k�lCy���B�kZ��RiΏ�;b )!��q\�� QI��k�,�4T�X��/l�?��s>�!�4)�2-���gF3 ��N�(MG鷳e�	��o��bwtȫ��:��w�ܶ&��.�i* p��cU��0v�.�ůd�25�m<o�
S�'�
Y���	|�A�"]��x( X��Ƌ��DN1��E�>��AƑw,[A�$d��9H�1\Eu+���@J����@��ULq~���!?M
�!_
f���� �T��GU��ƶ��R�����ܝB�8��%��P�*����R�|�k�}K�F�oy�FC��Y�J���TY�Ia������������ߨ<$hV�6�L�5$я��Y�m�4��n^���1x�y���u�� Wb������@�_�����W"q�w�0�D���%r�ٞ�G3ܽ7N_�!NxU��,~UD`�6N�����KR�iG���!��������:�}�J�)���[��3�1
~��J8��bfero\���xl������1�ōh�������J�&�y��A!]��D6_�qח�U���OGC��q��&��$R a�p���v�W78#(w���4s����!U�m��CDaӁ���@F,L��(y4�d��	��G�(�,��������[�:C���$M�ˡT

1���J�0� ��Y�RJ ]�9��(�V��to�F�)B�1���6z�|D����AI�`��+�і�D0��q1'�͌K��f�
�p�N����_�L���(�3	ĢV�X8�}�)(f]O��/�\?��{�@��E8P���M�(�*{��jj��F�ط���$��A����1K�PzY?D��qe+na�퉴٧��п��óF����}n|���z+n��������F��� ��>V �:3Z�bW��̰V�|���0��
͉�.Pػn�ؤ�n��/��d��BB��=��De壼����H+\�a\?]|�����`#I�Ch>�Ԁ��|���T���Wf�"f�X��+qS�.ݰ�P���O�[�iX�L��N?�������A��o���Kc��N�6����(�3$S]��H�*;uI�@Y(`��O�׿��/��/#��E�N����E�t�}b����i�% ����Tɓ��+�f�{v���9�ё,	�7/!#u
bxQ���֔������~C��h�Z�9���V��o�B��N�HQ�Nx�3N7�nc�Na:û-���"M^^�Tk]X�d� #:�Q?Dyl4`c����FB��7��U޽s3|V�)���F��H�ˬ���!�ɟu#�ŵk�N���dz��o�:�N���f0D�/<dG���B�X� �-�Я��xÃl��{υ5��4g- D_��,7�(n_��U]���Z�f�E;K[�3�_�+�"�c1�n�"q������� �m��#��y��ݜ�23����_h`���q����Q/F+�W����	�22�X3���҉\����wJMb���?;����C�J��
9[`�6ʤ+�h(����i�ri�<�W��jm�;���(W�h~]�'�#�P䷬��:MM��.z΀��Y 3��f�˄+�+f��')M B�2����ɘ�����x����3w���Ρk�렞K� �ˋOE	�a�j�D4;L��n��k�[&c<����ݸ�t��Qb�L��u�E�p�ҍ�r��̐����I����q)j��a�W�Aÿ���v��r{Jp1��:�8��̚�Z�^~)%Oĭs�Z#Ύ�g�=�D�>�duƇ;8#�w��T��];�$��:�h�$�u���I��Fڻ.dh����0صb�=�
 ������U}���	���T@&�'����s�Q�jږ�1I,��
�*Ɋv�����_��e�q�Ɏ� �J�uӀ(?a���&VO��q���[�q.A;uBX�ਊ�D�@t"�o�]L��;�AgL�-�Ih�J/]?%���r�J��w����q,M���y�QS�y��(�v��a8�z��5����t���Əj��6;h[�d+����8���c�#���Z`Ns��gI�umS�hm�1�� R4Ҭ��k����il7ېX��S.�n�z54�=Y��@p�hpe[sй��Ȗ��'�ޭ�='�0�Qi.��j�G��2���)fG:!��O��S�.r;���y�;���r��-,F��G��6A�����-�*{n&���4�@��]�(���s9���%J�.�1c��#�p�}+|���x���OV�m�|[R'�A�����Ⱥ���z�(�"�M�
�^6>����$hc_w2��N\��Hn�Y&��zcD6���Z��+3�����:i��)��pF��7��
�VZz0�r{xц��t�����x6��"��5{���]�cL�A@��d�Bۥ�'"v�O����#d�v���^".a��-<̋��/��$R��b&V�;H� �-fӀK`��MI`�x�5��J1����Y,lS���Y/�XG�ni����1 �ЖU�и��\z�Q)����O�\�8P�tt#�s~��0�����Jq(�m��0��L���4,;뇵%��#��F��:����M��à\v8���l�٫NN�2�^R��Ϋ�m�D�:� �́y��*��3x�� lGᖊ�L��[�4��$�;`#kǟS����e�C�$�OnJN��D�Ϊ񈂬\��iή	��U�Y��`�j��+�Đ�~;Q�o(��`DT��4�������9Y]A���&��:�SKCT�
���?t�k��4�KSBv�⸰~�#*P�TqC#�8ċ^�7R��]�<��Z�.�4Ժr! ,�2��.����\j���D�g^�M����`]��"��y:�Yp�E=�u�1DIE��@���>VP�g����}�7�v�5$C���~�k9��\��#P�M�խ���g�e�CZ-���CR�R��rvn�2[f���Z�(�G��⏻zy�N#N+v�(���p[ŝ>�L�`�����e��U�]H�Ǉ�Է��=������Za�R��;�㑚�af��g��E2��u=<ws�MoH��j/��2�-����h����s�P&�[�[�˟xh�T��B�� ��D�cIw`-K�`���q��c8��c��8X��ˇ�GZN	�W��i��5����f��5�B;�1��2S��͡^�=��v�z��DnW�((Q/�ڱ��~���2٪�C� �m;�;8=N-�����y��|=V2b�L�	yt���1WR�ҞQ���G�|C�8i��Ɏ�%���f���Ξ���Q\�8J]tj��� !P�9�z��s�ˌ���-6���z9������_�h��|�[����0����\�c9�T�ď�(*���g� <��sݘ�2��7���]Jp��� `LK���ѢE�&�<�%Z��LX=�� U����FīPw�n�MȪc�����*,�.���<�_���_EΔB$�~�t�ҙ�������G�m�@f�6=�F�2��ھR���œ�C��-�D����$��1+�`�:�u���O����5-n���Za����k�t��9�0R�^Uhe%�{�}>7� ͥ��N#��,����"���$��}fY��|�b��n�CS���� Z:p���#�����.*�
8�����@��Z$wUٵ�x�����Ur*>�8L���xy�����kڗ`�!��\���^e4ؗցv`U~��T�Tހ��c�%=nZ��EQ�Y���pD�$D��F��ml<|�WeS{([��P��UD���P(���GgUh`HvcK&C�6A�i�-���}��X�	��W'k�6��@�.�U�[h�Xjĉ��*M�ns�֕���7���XK�Ш���_.���e@�o����ψ+Е�2WK�`=E��g^�����9�#�ڥs9�-� ���6u(��	�1�#?병*]W��5���l<��ŕ�_�U-��/��ǲ��&U��	�,�&q �aO��f����o�Ϩ�x|�4�ȅ�SEo`�3��\�\�kKP�nSD��2�Bu�Lu���ұV��͘V�j�9�WTm���1�b��ӡ\>W�5����ܼ��J��c\N��i�
={����$�����������?����;��9F��r.�qZI�՟��t�ӭ�<}�|R*s�8�1_��o��4��{�c�V�l�u뿰=^���9Hx<!�[�CeF�t\�y�ҌT]�܎~-bl��m6�ѱ��_VC(���G��KP6�'�J�!����F�MJ��^g�W��J�6���LK��iH�R��~���9�9�g�y)݇ �H��(9$UK �DBw�Д�i��M�89NŽ��ga���s���De�)���3E�?����n=a%��$,'@���G�T�1S?m_��[���wBjT�e"E�����L}F��H���r2��~�Y՜J��/K�&N� ZV��	_�7�&7|u�<�A3_T��3��X�j���SJ�pa}���P�wYp��!�4�lQ+UG��G�K�4A��"���z�TÊ��t�ݝ�@�-7�"�S���dl{|��/�V�6Vw���%/��'	���j,)ft��_�Z�V�W�p%`FD��.U"�T�D�ݫB�i���E��f��l�ȸ�2�:�
5ܖ{ ���(^��Os3/'7�v�J�T/G�z(���Y��+�}4/޳(�9�^ʁ��ZO���h���0'�MьE.���
�2��Nx"χ��"ִ66q�0����Q�R?Ii�3\ddO�:AJ���?����:/���)�hG�ug'4g�b�u�LM�ԝW䛙 r��sK�5f$��!D����&'K�b�bRl�b�m���3c4����J�����E(o��R��n��e�S��Z�Z����S���:U��R�dn�*�<����1����FVL7H[�@9Z�G7U(y���N��@��l�����������o7/Jy�Jѐ�Qկr�J��ӡ���D*QI;�S����x5��N��.��&.��Օ,���&2�Y��&3�E�*���t����_��j�i�-PB��w���M��5�W�F��M@T�[ >�������Y1o���iҨw[OaXr�����*3E��)Å�����A�n�@��=``L�i�GGDg(q�ѹ)�Ĕ����u}�Ń�E����A�ѯR�YX�b��������(�|+�oV�41�Vk��p6a(kwO`=��|�[�+]Itq�q�yF�_�%�r/8A�Ɔ�9�*~���t���V��\)����Qc�V{<� v�$ۏ��&S� R�-6�x�_�P�:�铆2$�k���U���6%O,�E
�珆��'y8�h֢w�4��y�-k��jQ��!��o����Y����~hI�����ËK������8������_Z�Q*��#d�þ�Cm����ƫx���q��p0�~��&�̈́1^���������S~���Π�L�v2�(���ᘳ�r�Fj�r�B^x�/�����^�֜�_N���׌��$�X�_���_�H\�R����p5�Sg�.]
Q�ܦ�W"��R��ݵ�n�M>n�J���^�A�O�����V�@O{Ci�<��Wha��ꘖ_��+eh�&�[L��-˸��g�ȃW����o���Q�9M����Oy�MdA-BCN�U7E����*G����cC�@b�d�lN������k�����$<�����j��\�S"vVY�H�!�fR`5���S�b���NAlcQ��1�����C� �$_�%M�������iK6:��4��]>=Y.Z; ��q1���lhiR���R����$jK�j����+BemNn=����Ė����� ����5��ä�=�n�]���$��l^t�Q����4�;x���O+U�Mu�p�w21�+;T5ݢb��?�v�.!��;��,�WgN���Ջ���/���(�X6˿-�G���.�:�|Ge哨��DţhY�Zi�{���MN�U�F`kĆ,�~�x�,�"�?����-6�pFu�_MH!~�9������r=�P$�s��VR3��;���z;����O��~Rh�> -Q'k�����4�_�ckX��jg�f?���e��z�.��f�����NaN�����ا݆҇�3M�:X6�1��aio��I�"�M�gT!���8�F{N�2�k�o��[�_k�Z*�7\E7�[����,���҇�1o�������E��%lC�oRB�<����;�>?HW����%�����<ip\�	�v�ըG�/��gp�I�c�S�_�4/X���EŚ����S1 �u��w�,Fŉ�,ϔr(��W����x\Ge�ʦE���ȥilp�~����ptE����'��,���]͡���sɐa'�|A�;��	w���d�k)_�9 �����Q�U��zT�|3�c]E��k���ʒlk��ޝ���ۀ�~>�_ë[�t}
xz���5ɤxF��T�����E.~���֞7:��SG�l � �m��Bm��1�v�R.�ݯ-�[�㝬Տ}^�E���ei�9<� ����V��B&&*b��|�vQ�b����m_=��&'����3`N�Z������(qp��NCNy���|���2N��c�%3�4fM�[e6�Ӡ��X�y_���|����m��cGmb���â����K�3g�m&M���u0���V	�ԺD����t�^B4��m�`A�0;0�d�!C��- ����R�U�}-��=�:a9>�k���	& 9�Np���-a�0$�����=����# ��8j��WF �ʧ�r�;�˹����e?�(�IhE�Һ��Æ$8l0�t֖r��:��(�D	����8��7�@[4��eh6q�5*&�y{��u�%`���c���� ��/B���`)Cʢ��$�@��