// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
TUpNajgYo30ixWvuOSVTcmTUy+7e4GSKPGTSJcMn11UT3q8AH3gqQoasb61u/MF15YOlefg9wOtk
AOzm2cizs8FOSd6XUd0JKnxWssezGP7XaiNJ1asxa90iJjewh5LipmYeZbirfcWZ1355vzUT6aDt
lC4viY8P70rDTW15ew8xzEn2FFyDYaHPIpGq8pnoZgkynP8vj/YX+qZehyjTbhwe3MRKT62Dn7Qb
472FixDw/vmoVxHBzOOkuBTW232osok8q+E5f+P7eAwovhmVZp5Qrsla9VtqDNdbMVNJdV5pu+As
Pa0A1AkS9CxUfcMNBLSABXBH3eLj1ybWJ+ubXA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14912)
MhZCaIcCBIZjiUjpSsX83uheRli1XuGY8Faayeis8DgKzvT9Owc+zDijWrtnI8MpNlVa2TlQghKc
UystWh23Dl7h2ENqbeXLZzkMIAoeU4SM5dkgB44mlJbFs+X7dbs/TfPt34BPhB448qehPNrIHLN2
/2O2+X5wheYgmZfpvB4ymRwqG3z04evaiil7jCCAn+JFwlXkD7Lbh8lzipC5AGLXCDVcXizTdDbg
dRvv7uCct6rDFMvaaw+cMpIkpVveXzuVyDcS74CkvL4qD5Q8+Z9RdBLzCHQKwtyU0EAV2MsZDDXY
F/oLu3AIlhQIqmFLn2dGreqwnWsF1Hm0AtAV3pkutTioV6a9z4ll3Tc9FVEUMpJ87Qa02Z4SS6Zf
1CenF625MLOa+F4cbh8Df+RKsbrFMyxj3JfZndoPiwn++18zFGVMCcaxaBVBo8ttjiW442YVHum0
ABUMuxuN/lWtCvBvocs3ZdQJ53G2Ar734sSLv1gADzyWNpM7RL0g6g7WgufPhCRDDm+gZkjGXOfU
FHce1zApaUv8PLiE442QL8xCVM6rPI0pIO7IaEfT9y//1HlkSwgzHJ71zH1YsvfZmZ9v/aUnuGhZ
jki20xOJoYtQyGuqjMjLGx3hQQfQi1hJMqN4OK6rWuDt4U7Uepanbkdedb5D77EWL7IOt2WIV6us
s9UiCHSw4GvheTsx4geKkQJ4nKB5+1lp/gACn0G6KrlrI2/Q6srPvmHs8o0uchsHSzxwcXFnABDD
RuRh9Gvu6gRBUGNgX9UAFqh4EshNrvHl8wluEDhKQx5gpW4hB6TmLOLgTf4uuff457UFZ9ItyHUg
Eq6H2sVncGiMbYyxw8iGd4FhKY3BMdiU5ruOJpjKXWcApc7W8uFwak12b0LHiZNUYzQEzKoOLvub
rRfP0xiuLaCptnSSXM63kCQn9QKycN70yvahPdHsitUYZgwVfbPcL7n7JU2A3tuRDIR93W/LlMdp
7mLvRQOBxWrpOQUOMBQL5ehHyMs7GBo4uyRmBSDAxWMB9oWYHAeGYEgW52J4PDoAlxFT9K7D5Twe
ylAMYxWkj7ZMm7vLkEh5WBibXT+jQbUxTVwTf9b6mQ+rImmFhgPeU5p7qzqN5iD+0thQNKlNngYJ
AJ1f0TcKCIiDGGW8QtjfygL3TudClMmyAwIselWDpxVN+vgnXDGegTFblj02Jr2PaNsqaL4EQiYp
Bs3VozjnVkvNcz+8pKJa0KI9vhTJ/FnzfCbHZCsZTHD902w7g72tc3iBJNmy2cNypvYgVOyqyYZU
Y/03ik0ojOOKuV0ikhxNPY8dx0Gu+8kU5VCrCmkBuqIBI8FiP1JRG2Deo9lXnjELgriUeKMbT/y0
wFQUTR8Ayy1EIA+wBn3vszOS+4mNx+ZFj6iljQU1xKhht+y8tHuvJQ6XHckPvWTI/0KJBomWCt+4
wNmQESRVLv/jxUlAlkxDlzm3EDz/mXVgnd1bfbaRYmCi2Le5ryCo81bfMU5VBvhrTqmWEZmz6gIO
N6G7wXr9d4RcwOkKkvfnI8hOmdcY7o19L6cmpuzZij5/r0rjkEvMsWA+JGHatyQ5K0+xRQB2q5fe
iUvuNGxnZHG+RsY1fwarCXHsYwB+Iti/g9MpfLe0+OYFdxRZbkWIWRnNEMZY6vHTcJbvT1EF8xbh
tJEE82PncNYoOl/VzgP/j4pa3j4aDRhTzcnhtKFcQrV3Oh7ytd476d3+Tk+twKAf0RXA+dHDWnCe
RG90zbdJ1E7MllFHZqtSbXTLCiJpSotS0uPCsnrmXD4YlN9SGt1uieJtzJsmmmixhYSUvnRll3kC
fX8AUP9P9tujCsPpQYluzp+cgt0CVT3NsAPYjSZaYA3JBJKmRcWDAmEGgLosBOHeKSjfGA0tsaF2
e1lPzSv4RvYzkTNr4o3XsEfzg/2RUJnSg5Cw8pDS3N4An3UqWtdrWj98Pow40ACtWnEiauU+m/+M
sUollZm6etIgnrGHImd1RQ5A2jdKagGi/0i9JeUbp77kBMwiyYEQn/kuzuSSzYWFBjxKQWAn8fKI
1PEwY2BdVlHwAz1Hj2U78G2QaVOslAGoCUpgfm1N/Pzgy1d1YkkRV0C6TifHuJBYKMQx/jLWUnyT
2KC3SqjgXV4gXDhKVeVgyQw2lkkFmriTsL9ybSTGFZKX6NJnYJngkY6MmpUdKlUZRg67BqgofVVR
pTKXG5xBLvJE9FB7FM2w87JX4NsyW9UtYCZhP9M/8D1AG5tDcJLearqSRgJSX5U7PiX2yeOaNLBJ
W0ZM6xOV8U6njSVuIW7gXSYEYm8OWOmiw8OUeP6vpXqhLoTtV4kWxn3BlhZZpFLzE65MJEydTyvo
kg52ojCwFa7DgvPkRbYXmKwQqm02Vgr6lzZaVfkQEvSnkoMh5RQ8dBM6ji3WTJdIB8YTa2rkwyL1
Est9T8thYRXpggDFSJQz0x8d7b4U+RQtNQCkKf6BAr6ETGCCYQgSkOd3hlLwy/EcoxXkTz/v0wqO
fW8vjnJzl741eAHHOTC77D/vuHeewXUU0n4Jhwfqt3oIEu3Nk5cankYU7CE5tzjOtlf9Yc/LWSXj
MapTQlcuOSHYsgTo2EsFBMGjUvpjDtT3LjyliprzuLy4DaFSNDLo/Kcv/A91PMlBQqaUyywZfMQg
MsQd7gyhOWYpsE8KPglzk4ART8EOnMvDzI3EZl/XZFgLhsBSvtYED7a5ESVsfIdIElaMCHv4Zxvn
UQt9L+GeK0xGxWGDbKIBa63Fo6DJg33uKTQ9o2uEQkWpULVAl/8Y2TZ2t4nXWB1QSlm2NelK/cE0
XfrGQOLYtNm5rmmiOC6OJtMEuiMqJ0EIFJ1eoiG9w7p2b5xRtqCdq8MiFpKE2rBHfj2FA58qWo5q
FUp8ASkBb1eE4t3Du2FjEoYyLA01KAO+d+B0zCMq+aQ8GqkIl0k1WdgquUKv2qob8xu09dtnEiKt
Jx/HFjJphgCgHhsy+ZRPerFLyHhzu3GJ2gmwDiH+OaVcSqsc3JVyJtjwKZrpAEzAjYVDZZY3Uc2A
KA3k+ke9koNPNo0M5MhpXlqEU2qPpKxEmx+oddX/PGexwLaWOUFc2LSNgBVOt6GjzXm9UlBNFeUd
exB46hvlvWwEQdftUtRnsSPZrAbWVvRZEOD+X6vsGMpKsBGD04zwPSW6L9oGdG2skjODznB7WrG3
rzYRpyla5INDOPqvNEECdww7YQRz47Y4mnCxUYkQWdraQsgWRyOWwTtYpNI3bKCluPdWQUgGlEpQ
oklI2muOd8Nki1XoLJlrZt2pPQxIQCfxnwlbXQaCDboDbNlr20VMwdKBaqvMAp2o1TRtf5T36Fkc
lEsQMMlyB8DyNPLD4u/fqsyr/4garH+knUnRBUnZbU5X2upvhyB3oTjBQP90p+8GSmNR/Asa0oMG
+7AbXQlExXzHiC0R2VZHlaMPrBS9812L8h2Gzh/39QVqzQvirP7LwgeCV5KeTT5dMA0G9W8IAU0+
D8sFqwO6XZssqL+ltSkLC9TbO82eGI4TeOT83e6uTsyM7y2lYkIc94UhwR8phd5fZG8vBPgFqrr1
DTv+SkPoc3yDcdS6ZVm7QqTUMjvHn7DSn1/PzOmeMzT+Xwa4DALWRP93sbkicWixoIyQHXQHAkUX
Irqzu1+0fWC+ueYno8ix8FOgTPuwXY6W0Ki7/ObP/mW0/7IBarVb6ylWLV6LjOc5oHKiqGwXLHvu
V8opayBTcmJBphKvmfLmakLjcAbVTHpyE1KF184d9iQVnS0uoXTF9boupbYT46dqL+/iOpNAQXoQ
KagrGzw4sJgPZ0Il0aWYz0rnrKl2uI/GdgDWGF97Hmte/FkaMHgwYsMR4fjCvyPMg52diJ8QhwQy
D5f6utQz5AJqEOs6meO035HFIrctWV7UCba7UmZHlEsPuQhKV1X+AQhouBNx75s3hgs2dpzAsYku
pNHVLNoSuF0Vt+n0LUKWsPLmTHsSLXaAAZH4eR7jCBqcx9oiIG7ndHL6DNHLp0dDLZtg0NHDM4ck
zP353te0VSYcwdfPNYO075U90S8nEJRIacrJEKeLXt1tsx8aeU3jQcJvdxxI3E1pfDlAWMOcqwQq
IygzfBb6opzfRDoOOsUx7I7Cw6n38wwPNLLo40Uu1lo2uWIehKX445Sqcs078Qq5hk084lTc8l+D
gv/eq7d4zvG7UCUHMvpVIgz+yKdxNbJqhIkgXY95IimoQkjdnviOHPBAeNj68iWTHRsyRrcgheLM
Nbs7mllhMMwSGdrNWe0A6himS6qx0fSTq3jzXGmhzsgTTpVhURk+R2yVJhKosiKPt2UfKadHw1P1
1s5zzYDsyutfibDOgEbOWkGoh/lEdm8tY9zxBo2bL7fFik36WNngMFcQk8YAfk2dJzqXupMuxs2J
1jUgVO8IlZyoOpLYEy2+WX+NN6Bt8XOkgW8TCrBiq7f+7h0NNC+cXmJSnfh8EL8PTOboO5yvoOU1
8ykK+1sOF5PPj049JKhh5vUlUuhbfTio31Et4ZmNo/VZ6CgkWa9Crw5Gaalm6oblqHnFWklCB/sG
kJmlZ36pDnwnywP1PNJpATEYKwuFL6qBMSNoI7Ba6sI8fsaDYzcDNO0pQXu+vQfOR6Dq41bqS6qT
PF/RpVzRqvkQ1mtlaA4UPWmWhcQbFpHsl/OGjuXLAnyuZb9jnpicxxA3nDBbay37YdJ+wUY95lBr
SgbL+CRnNG3HfQw37XfNfZ6rdiCYkYfODlT2F2G+1tyMUbX9sTaXcpHl69vkN5GJT1mWvjTHQdMH
LBhIrmXSa+9uDzxJ9mVxSJlVoHh+7BYZtsfWI90IjIucXIIHLCAqihrJBRzl8ezKWbz0RBuLljdK
Gj1CvY09bqu5c7sb3TYDJSR9JtCYONxJC7R5AKUeQEuX3ioQ5FR1zwVRdLmfD6IAhhQ5k8alxQQF
TuQtwMVM8GhuzyNoTLeU4FBAXa4dsGYYjoSlwu9wQsaZPyCaXoZVeRZUazuKlZr9sUAYbCOXLRmW
lH8x3BYEU1h8Asg1+xn0AnJQ/g5R0v4jr9lWAUXN5UjGHwGbWbRuukDPDW6+mab8paaHTyBg4tY/
pVpa4wOH+SrlqVl6V21KhXL9ZWw85QPUzAH8PCHhkGKLux/2/bibuGK4+HY75/6vP3OIM8OX1EZw
KMEZwxD+jxP+dtait1guvTf/i7aB1JSue/QCM7IXxvzpoOmelDjSgOo/4y9E+2wMVotvoa7ytFn/
0PmAQ69DpiCy6F71Hm8WVseVqqH/sHR08o1ETWqPPumYPAmCroM/9fPc2QlHsEZHA0644DznZgxz
na32RP+S2t204fLAYTGtL8ksOCyw9P9qRx3HQO/nGmT8mnqW45EwHW+eOs+3Qf2qUz8NR0KBfDM/
+NqE+y895d79wL9sUTWt1s89qEuwxD/E/Dc1ABL7DlzEX47wZteFr6DrNLhqzWqxY4lPmNQHPsHM
ZlRyOmp55rNrR4a/66tySHZ+YhRi0rqgwDLkezyK6W7/QumQWpWX/aX9hPShMeSzwhnqTPj4axMH
/yYrjdeUa1fdx1GMNF9e3hafaO8kR5ct6ZPuXSdGGoJfoiVDf/Ca5665uVxDoa2/TYQqGYhLSEGG
9EpeFQWgjfQ3puTxi0r5HMApwExY6GLhnFuo2pCmm8T2G0VADSXANSR8GdySJOG7Z+2uV8bmctXY
OGcLaDHF843X0PQwdzMbblx3Q0axDFPmmvC4wCWFYhgsfsqyc9L4YxuckwOIedF3rTuMBm8Z1FJk
SRxeY1TBb9dvslVzNO92Jd5HJG1OmDeW3dgNNlN9mKsKjb4jxaHEKD4vy8wIoRJPMzocfgLK96bi
wM4c1RlyRRL4o5UtJXZXLZ+B1PH9LkLq6RImRahQOL4LXpf4145nK7/E6y2h9MnyWsT4jwZudhSM
R1nNwuk1IKQIGnnibfZXguO6uM6nYL/6a2Bt8dT6+GWWyzpS7kvVX06/OMEcE3ekRtsy+q/Opdxn
73t4AoXkdKTa4JI8XTzFJXHiWUPIKHkRamRY7l/jbo8AOFYof6SQJQrnJG7Pdct9FPD/nwyhb+VT
eATGM7HdDjBU0KUzItgJfhKu8S1YUF/AXg/4pYqmou2oCWzHYLEpHsbx19zniabeYqPg3fwp2rU/
gaZpN9lQ7qFZifa3ibINA/pnlQMWAcRWcKaqEXUMDWcqX7+GZ2UOHeFQmTzNYSMVT8ZQPvf7QPyP
wErTItGL/U1SuiqWoKCTBxUvO6UHtAjyhdfVgJMkj0CY9OYNmYF6Ai1gY64UQW1YT2krMF3n9X0X
AApQu919680qj+mg9aquiPP7Hm/VHdWB+cOa7gVIfCOsTKHPi2hn5ukOvEiSfVu4fvQjlEk4BLBS
YslYRzpLXj8Xf4pzAdhrOmEVDy0XDrPL8M31Tq+KFNRL3jLdAMGXaddqPOi9fAapE9HrtSgQMno8
7Wwe6vMdAI3SsxxjzBSC2fec7TQqe4G3nezPM2Mc8jOpOLD6cumMzJDdi3QYOZAJcZGh0u1ho++S
kLXqlAUKkE5aK/QrcLWPDXT+QxaDZsn2mLdymy0WTrV1ryZxT0D731ARwZi09dDjGVzbQo0EsrLq
vUbZp9REKladw79y+LtfBb1ovzFV2uVj6Een1eXGwwFIwimSwNMsRF18DbX8MORuHsqqn9dVEjhd
JGcDTRGqPsyTuOaiRe/Lln4mGnXH0WfWdL+Y4cNyDksI98GhV50SQG7LDmItzmFCEWJBJ2MKTCrN
r+dgZy5iqnccSRUNS+XHhuNlRx6CK3xZpr/JzGzIGH1CNnmX1vGUJ8jMy8CxXKzhux5mLj03rDwg
x+BRs22vBLc4rXnOxVuryvaNql2h2+/qRzyr8UJyxvCMo3m06FKGDAy5eAxDxzm+OiDMcAv2/OGV
moy8MPI18BzBo+M/nfayJCkV87BpVWRv3JxpOs+z90Zjl8Pt0OjTaA/veljmhEHeE0rxrbQ9tAs2
XEBrglo3JTKTF/DzDamvRrFNpgZo/VmQhnEKEyEltrrV/7z1u03J5lf0dq4Itv6kyqMwYAYlnzSW
ZQ4Vh5sUyxUGiv3IMWlfFci5D8eXQWmaKV+15/oUOnzfY7jT3E9+0zDfiGZSoldijj1yd/nHRU7z
SyXchpnMo0tlYNu2Hi5J3Bz/PZll1R0B1QRgMgyM8YHKj+4g+a5lvr4aefZvddP0NLBI4mvGb08p
+qCzk3s1Z8hAhY5V37+wxTTEOyW9sjz9MJZ7ORvSL6GwjJX10hQvamdZFj5JDtsC3WVaNn4712Ty
In0dBbFiaOQtLoTV29pwwGvDk0HxOGBDyzvGUDxH14y2CNPkc0KdfsdL9e14M5TptrH69EagiY/P
4udV0qQq/VcuS10pCn0A6efZ/i31lDqjy4QYN55bDkhWSRsPA7cjptwwkRoh26e08aIl8J71SAwl
qhOGfwBvg7iAMA1HSN9cMQ1kL5Oh7IUclAYsenu2lVm76WC5z8Y3Yxqma0MlJDcrxa8EtcCRWs3p
bnRpbezhBpXratN50a+aAquiwlyyT68QRYuL5BA7+iU3auQ/OabJCi8DKY/FoEbyqRSnxGBBdzme
PQPRQmyh4apsn1Z1xZvsiPU5pE5ZdI7cZXsZnnlJqO0E8gmVRsS3T9mtlVI113ff4/kjYaXHJNxD
FbASXriLleYqMrAynLFbEg3j1IyX70C/KHWYXrVWS1U/doxnFLOP9KkTPkyg+Lq+qGAFV30/ZlVb
OKtJ8ICUhQKU9D2e9P7TZe8lQb85fzPWoWDNTAt4cyaFYeqjKQbxfcgknnInldNpB3aY1/dwPVzO
vOuj3ccbtXjcrk+1/6Bw/fH5aJwE4uH2bP5ZeIluu46svNPniH32bESJrVytKIe5AE6JFma35PcC
/hd6WTuv9Rr2d2mVHtap7eSWrZKWT/z25uNeJogrKNykumUWjhz5scixmI//55ZTbnlXdCp/7xtx
QIwbMj4u6eRF912l6dnqmSouGa2MmK1K5yocn/cusG+D0hUhR9RY7te/8ep7avF5iLa5PF6Wxb+f
kCq1tSZGgBNTkFEhaTtopPl49UHmujE3EZz8FzTRPz2hCqWjH5SXT5bSAerBAGQ8cTK6Jrrm4hLY
bPZRgJmsv4BFifATiXb9LAsHsC8B+aPXUkKwNhvHGxt9xyKXHbMp0asxX46b9zgIp8pz6flfUxf/
Up0h1HGH7YfiGKSLK1kvqoUMLb0jx0RtEAy4PAqa3oqMnCgjpV/nGI+KhFEbLBt2NpAWwudapVVc
pmF25SxErTfefeuCKp7B02j+MzG5M9nlHpk1qlFBP8z72WCraxuWVwzzxVPge3lnl71nNE9nVDYO
McN8+C7eNumAcdsgAfP5FXk56LY0ASPu5tkGJpHrbmGQHVcq2fD5JEIY9in9/P/3gZab6J5D4DHc
PuMJYrnqfPoonSO/GRlK+eBM5G6cr72lKA46mal0XLQrU+YwZD/Oyv2ZINs35B06uICIHDouPH5T
UIiQ4xaw4JbgE3wMNl7gXwD62MTW8Ps7QcKfDX8BZG081mMqsprvCP8QjGZpgpgT1p2uTOZeJZ4S
sPN0g3A427lhZMZyzMpnBFt8gL7RDvDA8/7rOXoRvxBES0waqE34xg1gajEdzcPUEVm+thNvxikN
n2ptX5IP3q0pBkNUvcMUWCM2r0z8MdHhHFgGfq5DVOk/cpqqsQRjmFIAIs57GgPkO721vdVNijzJ
FB5NAELWrgn6NdMrc6xOnvk9ZuhLQQIledVW789TTsL+CEFxW/BbGiMCqhaxTcINATtMh4Lwxb4e
5oKB3IMM1kVvm98bwB/vje7p9WDDaOP6rnBhfdN0O9Gavj8yHradj9Ts3u2fww9qV7ivMdxOTF1O
/+LNA7GGMiY7g+2URpawW43/3BNEbLcXiSsn5gmkywnchd+KqwPdRZBo8sgEhgZcgM3ZK2ppfDuM
9s1HUii1bIoZ0Qi2AWXVxoa5LgmzGPjp1eVIlzvt1wKiLIh6CRKH5P7vX2kFTaj688rIOtvaGfrR
WY5cn4IYkI42cQiyY/7YryPlAtB1CZYfJI7XnQDb+F17I/vW45CRezlEAc1QCGkqBDqiSpUpsKro
o9LFaz9LeXBv8LqitdlfJBTXcgtpjL9+H/0z8l1KRtveiOLmdChJfKnQP7qAQQCy0leoS8IdeQBu
aFXWtvgVRuW41yJ6sdTbHFF4NLOKI9qPC7iRST7LEK6eknf5s7SLaae5JtSG4cxrkhCUc1LBPFd1
V2K3H2YAcs2qUNZTImb6gvu+KG/OADQ5ReRJ/sgrKZUIDEMW2qSQMo7owxwuVKgJQVpmEba2blEL
xeFdAT7KM0isxecEgyJyQTSYQ8gwxsXx6yeXHja+oEllbGjonGGFO/+BwRc7yHjZRHRo87GMbBjv
RFlQ/fiU8t3Pnb92avh0EUGE+UoUW8Y6wYh1UK98V4MjzU/vKrGy31Enxpyk9iKAgRD8+FNvw6Vd
sG4kRW7XoBYEiYuDhrQ3fC+EVo/7dEU8MoVV+n6zK8FMnlLGNaQ9PxHWVWrNola2S3F30VVZQcxU
fxLeQ/omHg2ZKlJyxSHnAJDxtczxhbrr4Zdz3CDJorSRp4a+qaUo63lkoQypdn+INjen4h0huFMv
UDKiWYNqcB36WKOcoK8mvCuGoONbdoSQGgYPkHA0cnmeOytEyhkxxcDl/+GaN9SCZCXbDDfrj+Yw
NAzMvWZVQM7Mmr5EjbdbWou+mCzHjRQ3tNC4uPIyVyrA3RspSDbCCW7kxf/VGmUbfbIf3u+OGres
gtDjmsgyqbSPDLdDzkRM0ZO8OCSIJgLn4BA5+toM0hd6P0E3J4F5CDR3mDoYAeuUgiLKGz592rNW
vK1o/dzgL5wP709ZX7qA1hms4qYFrhwFlr4JLha6aCdfSJuIY4R8WA7QL1njznD75M+XxKmxvNcN
TqILP6V8dxBU4TtD4gXdch97IBxIxmlqgrefvz+wVoDfOY1HZElZN75yHmMHnZy6eRW3Gv2AFyZN
A26WwotGUOWeKYVDoLtiwloudAYSHyOs3a0R670CgQ0tl3TJg2+vsAuFtJ2rD0qc2XvQxm25DreA
WEK3PFVW+m/3OBdaJfI/0wyDss3EQYvUpK2ZqpKtGVK/GONw3bROMBJnUVJ3KNlQi4IZ1bNjHg26
jOsQMBi2Re+qHJZNWdo5Bp2vdygqC0/zxC109PGH+a6Bl91WJQDwW/T6kofPO5eTt3gHYmBcs4vc
80fVMmg5gs6qsO68sVMXvlsCL6u9xjhvByMckuptjnogsMPpxwZ8Tn2bUjFpRSmwAzJKmziJ94Or
I3bCXM59PhVVAEqAYtdihAgQWa7aJkzNXDQfZuKeZNCgSwjtAWH5m+d7UZR/cu9jfGmUBmRQPGj6
hq7RBSCoKSt+UfnnEkXHNHLqdVpdMSNV5YDBtHu0ID2DNWz+4eFGQeV6ymBtNiUsOZxKs+AGQiYG
+lAtUXWrDfKbijFBby4iaopftq4blo+/sOERm+4BYltMH3VmsfGP+0+0TNg8cjbB3g40ynHZd9YU
5WEU37p/NxYi0DrTcrIqWxPioQJzdwc/zjluXJhbTiKrPT0j5vhlENoZD2P3+y75CwUqV/aIUYVP
XrdUbKYyAojEWQvpaq1VnhSfnofA4CW6pgL0IqKf6hR2hNMYyphq05jlGWdHG+rcOXFaRJGZs8Ym
aOjwLl0awr9Ak6nclol/YUmcmO6uMmpnJtdqhQBSfC78Y3D9ZMSVffl2CcfsSk7BS4ehzqriicw2
C++ttZKZh4AWaLdDObaU7Xfy1i1lCO5Aqp8s07w6ONbW/qGoARpzK5tRjQbncLIht1rr6NIed/rH
WtIzauALI5T7+6OQE4bpW334bVgSgxN7mBIjvIyD057uc2SA/g7MUuaqfoyZVoFTtvy5YdcGdIYY
e0sca9nDqqocstlDEz3dY4zBDikLsGiMwd82x24ofaBIoiMcHDiu86kLbEAWkx2Nh6R+D/m/0vDf
MYIPCYO/x96NVjbwKskFXfFd0ArhRUcdrRzWNtIbtOI/DkLih228yKQvLa/mOCJH8j2/2tsFi7Fr
xHB+kitVPcngJRwg8HCWDEkDvkWpjBrQoUSVsZa2wwJOZj+4/Oqznq/kP8OYfnnvk9CO5uI3jlKO
MgM0SIo1oiyyKCk2wnOSDvg/qyEcXg8mO16zpnPzKIY6KCEeDnwIrZ4uGXLF1PF7KncJ0g5gxi5i
SvTRam34fyGm5zCw7XD4n2j3dwdMl+LzRHr1USLMa5m+N73uF+xLX9YoVbiQVRteWODz7FvmtOwR
z9lJAJRHmH6OUAAtjxL1C7ALkUh5HGiDc1E9ITJW+WPBl5mpHji19t5bCWZduhXWXdsoW8TPQ+Ax
hliY8UAoDjAZx4Qh6lsrmpNd3g4Dp9Mc/xaUYgpZTYDak/zpF0uA19zq9f33J2Vo/6JW4mMUFR6P
YGlXjZj5bsF0ptwla9cqdVDh0JgJ0T5Czr9H8c8p4G8lbujuYnBO23L6F3/35WraZ0q4ZRKLDQ2/
OMTmRPyKCeWZeE5ONL+3YgDNMOP+REwRU5Y7Y9zFDiRL/kl+/M2Eq9jMFMXCKFpXcNXQNO0TskO7
Pv0K7dheaB2snOOoqep41SNF9QWrOzqQe66EPWfLbUek1Nr+HD0Ksi9NOsN95oDZrp9a3VMB4Pad
KyR4SALp/WaHEgHPnu5HZcLMrXMD3o+yG+XRtQaI2qveOSKtrYJaBXDO67XUairUXEfcXQCA9dR5
t3yumlkTbAuxARl8/hQpDPQoFGe5p7j5yym/QETs2qyga80pPDqsgCPHaI90X/3IAuBhecEV0pEH
nKCH7TFNPyVuezTbfnpmXCG2wCN8tB1fJjboQRFJ//2dZbBPFieFyPsCGiivX4b94J3NYT4Opl5Y
+GsQ2G+NKsHeKy7yMVjFvJ3/Y/HfUaLfh/mmTJ+sXoTtq9k+/HD6IUFToPVbMewdVNTnqSVJZGQR
UCMMEbyZMuoHhFEQh9S18/TIYoVuWV4L6W6y1Kuh8r+VWUFEY9/cPyAlitMQfzi85mjDre5wi5f9
hEWK1/6xo9j7WwCzoL/+1yGJxrumCRrTGRp6f/w/phlq4/YFk1q5+7EV2MrIaMvSsXJhZqAfqY7A
RywuLMBVq5Wd+4hFPHKS2eGrxPru8AgpRAI7E/XNbbLi+KOfWfFleQU92H7CXS3wVyWV+OLPT5a0
bPZWUEx3L/pyN7QFU5Ke+uyDK8MevzmxBodvMBbV4SvhfjR+6jefkhLbs9m/5Rl5ddKdnWSNdpsr
1eW0Dowkl1NV+VLzcpzuirNNWtzGbMJNeo0ysLaxSUh9q0v/cyRlNfIkanDGCpd2KaInwzDwYYXj
XhswZ/TnKran8PFAp0V4ULApE/wU3dJeRTdga0kbIAH6prD1uRCKtqsITRtDWv0zGVHJUfvYs4v4
rQ7KGMGgTFnH2hN65UMIpxeZ77DOp7ySbxU9B0nkbfcNWBCJ/MG4Pl/2hKdvxXr0RazSMn1gSclL
bTexIMyEEquQ/xrjVY/P7jYul7oojdqB1qyuwiuoSOTTzs5mQhhy+ije5kjr4l2NvyHrfsyAdS9z
WCLN8tFu05gbNCdnRc/oVm6E1JnSrPjgOVxeUPlYXRV+rv75+4B/Y2aV4OItd5HOUOP0eNv8LPM1
Y+rMIXO8aIv1mT5/tkudHvDaoKNNfkiVPbQRLGD7o43Fm1MYi3tahfxRbRT3jNxzD+rmBqPs0isb
W9/FRIWa9eRJwjJcaOBHoxDCplFg00w8omrya6bjbYvYlmt6wfjs1Mbg2jWtr7rZZuidebqkEWAZ
IBTXDTWkpJVjm8TXynyyQ3ivGb1Q27klEqy998IsegIl3ayj208uDa/2NcI1I6oie78WGA5bbvkt
d6YEOq1ukLbVqS2OsXQAMLovlcnmDW8NoH06kPUBf4/cSmpyAIQ/v4/V1u3L1TjQveOiyk+5fXBV
rDmJt9+jUppFqogcTnERBYzZsxQ/1quQN/wJxWOv64pG2qMsZST5ak4pHeKFgxklhhgQyPLmvkae
NtrjnM9Hjh3/cR+CLwGWE/5v9Bc+0Wm17Oxciw50UYKJFV+MgW7Xz+5yZ3cIY0W7DO8yjvpj/Fuc
KaLMM29NWpkuP8+3tB8nocccsqigYslI3p0s5ZZUYVnxR1aug5dN/hDGvkRF0z5bwv1FxiUOPRZO
7hXm2PIkZAPHH2VK2d3hV6Obwv6UWMOezuk8QIcpQb9sbvv0zOrak4bWaPgClpANsTaB3qQzWqVT
kbKyPQwlSbAHi+Nqqo1Z21PbuZFt/J/XjG9GpTDPsat5eFvp7y/P2/0FtQtLBwujEBSRj35CkBuf
ofezXZ+JYx4RG+07xOSobDv8PpakIN6X70uiuKgn6yC8z0IFAuMUa96v2GIrzY5ytH+u+RSCIwJM
9ha8FTinQ/nKreRw6+ILWkbwE+sJmOv1ybO8dsSEtJCAZfZtmmwvgyRZr3TrQsRQUlvtDHiafSId
Gd0xKfEJjiJoeFSgAY7bYHasat0EOA0P5TuAmP806+nD2VRrLSM8Wcc5KUC7wLOEPpiIBsBDCsor
95WQh/Q7zrn/0gk1r43T0e+bSIYW4LRnQ05uUggUjFRUSLTq/1eMiZfhILkLUjBmkfzPqBL/yp0V
wgHhAAKgTNT4vwUpsXpThXG5nNhU16xftUhv4SpcP+r0bOzBDRorq7GdRYhNcUf3w71aEGNVqb/4
9+0IpYlVpjp5EzI/JlrS8aVE+w0dEfdMFNq5DWOKdk/ObyXgFJ7P0fSrN7A5E+a4N1NYDTG2XlVD
qQQpcqRKDqk7vK5q+QAQNzVS/pMXHdVZyXNpzFc4XZL+jGVHWs/WW1h3CaNVnFiypzLWW72OoVE+
Ea31MwX7zXxHx+jR3jZz5Il8JDRsG9hG34eV8DzrNAi+dviHsPI2R5ZtoT4J2CyVNmi9J8IRjvdH
JoC9QoMJE2fnl44yeUjkqv7SVz3zyVVHf3Bgv8nFrXTXJqcS/ThKAetQyBPb+XB128HZWJEA35HB
aMg9VeImHAJg+2pj+Ttj0jQoaBsx9D/+37VsfjmCR1yZUURr81bqRF1ZenFuaX872veNit+NpA7W
fBVGetIEkkOy8KAdHE9wNCw1rOMWhkAkLjURSDeM6/3aifOVKIMtdmQBLzHBDFMIvTuaymWhz4pS
eq2R51BFSb2SXAIDu3MbTtgL++M69F1SQWYqtr8AWIsLkN4kr95aWUXkiroso+BJLsSdzaje9grn
Vzzfny+JHb14aZY50XdMVHuQViXdRWsoJ362RShWOiS3wutUkBfNvG1yhOWR9vjYBqor4FxHAHBy
wryxnRed3qhwLNOBJASiru8DaGa4HYbDvvfzSWjNwRjZwsaDAbp0u8m77PGJRMM4K4FhwFXDcVeu
nVctMzVn/f5h4rUnYI+DB6geulCd2pIp5SKoil6/ySFnh8U6PfdUSlGlKZu+/7a4DZ/l/jdjJ4ns
Ne1tSIwdrdxwxBH6A1sVYGZIOwNczYK4Do8PIt6qCml74bJqgw7MP67e0MyQBB3MEwJyE1acIA4S
7D7lcutgIsX79j3cQS6S0OfHGJoIJtfAZpcghVAb0gDLI+7Mer9HoExmmVhhp3prgPc1l1DM+Gz7
QdGuwqecyxOksg4+741RPYaeRsTwPST8nlcPIQyTEkjZnFBJNvSqHIOl6Y12Quz0yoUdJa2mwlv/
sdye/twcrjA1y6bkg+Ue+dQ58Wq247pAFd6pj9O7ejKPHcrZaVuYl+c1mcZ95Bvjr0z8Riutsq/W
wU6mktGOvS+T/QGZUyc71qdr0gDJSswcIvyOQWwi1a7G0Hpz7B6fbUT81R5yjy3LkbXZY9d0M502
aGKsuNSj7fCjqmyBCrLBxo5nTjaO0Yx6epvvIs9+q6jqJ/FRPRgLRzeNrLtPipIsm7X/krkGo2+2
ZhwGnI6+6KpKaWGZVphcMXu0d2zeKTNkOX9Ix36jXOKGKwnrXOZ4io3K3KSY6VCbj72Y/03HGshv
3ISGMZdT6OTUV3cieqF6bCR8vHedF9/9AMMwdq9ySsZV44/4Tba6IzSLjDp3CCE3ogCr0WZkjbda
2NDhUjUwbUSJw6Phn0L6z+cx3DSO79gDkQd5j979nRTMXrF4f4uKuVZPWzC1zxeDlm5YBCdgpDzf
R4tzC+JKQ2pPcnYgfV6ASU6A64PkSvSdDwdfltJWpSbGQ8IBw9Ck8s9RJu5Yq8C01tT4LRaJTs9Y
6bl0Foqn7YWwa43wOJs+W4KuruSXacmkergyUP8I7td5T/oTRbilGuV8DC5uLedL6C2Kkij3jHwD
lh5lXtYT0zNIlNtWXEnFjLW5YcPo/m+OeOSRhNFuLY9yN+hh67CBPdPxEIzTIXEtezuGJp/cWR+D
KEGPjKk5wowXCV6m6XxDtJLqnR4JZGv2z8hTK4rdgSbBoH59mxJopvOcYkEPcHlplJ9FTtnPH8iC
9RHrOnUVNmup3b5/yU4UGPsRNrquAtgua4dEgEazei/a/zMIeU7rVc/KXnN6xOEIA8t/mGFKlXUt
OTXH09aZifRWDeEGE1qBUMlCq1Um+7RRf+v6eYOll9ZRhx7IUd6FnsLtTPQZK6cw+l1T0+z7fPjb
4l4DeVp3DP5o/Q7EQUgsWvZ1MnaWV03sB1dKmq1urspoVcCvjMTwUD9FQo3LpPvLlHMDBXiR0RfF
3j1sJdxX8lAZ5hRtoa2DABF13tNpY1xC8ry4hniBCD8xgc20v/Jq0Q56tHtEv02+POnT4BzGzRaW
4wqXH8uJJ4k1EOaTzCfb0rr/7y9MI++s4X4uMIgFUP5LPsum1j0tSBRRn60jLW5OWRh/DUWvYUYe
l8gd4nKApi51BAAl1mSDo0qVI7mZpTJWN5KiexbhZ0zqzwDsv0staDt2mwKkLptZDGTKlrRVLkTM
LoMV8H8GYByIt9y2XXXftJcaiJkixypkHbwgSmKJVIGSx2DVZeYkRHRyV6qT+3IHzTrueytSlKoW
RHWRQ+ys3/hPdQKnyenXrMfZcwTR7cG0H+dV2PpasBPq1j4ww+XuYRzJzou4hv+QaHb3DDfw530m
PvsVSsjGqIVoYXpicz4k5kdKMrcE/ci73HoJ4RDtYAGRV05FfDvkMOxESuFjPVd/iM3Y128P1eVh
3wxB9L0+OvYHK5dSHkwJnid3SR2VqMAX2M+hRLBdo6oa1W3KJ8Lepb2wLsFYtmEu2yNyItzZNAZ9
ev80kxEe3yO6McD1og6z3PNAbRobmbJXoNAS4pt2Dh+pYJCurrrnh9WNC7nI9SzdnLRHc/yAuR4C
T/ql88sptyNi6PY3QA6++tH1mrnXri4X5cjUPkVBhfFELSuu9VpWXF2t43wQqf3zgj6gofAver0t
9bgztI95Sb+L5KsyWAX5yi+d9O6DkUMI9a0/ya1XJnrr/t5ypQWjikEEZlb59pgndc2/LrTAozAn
JlElOHgXBlhMBRHksZSlJ7jZe71hEGc/HI3K9T84HhGDavag5PrlxRBC2x1iMKrRRPUVaYfNbo0L
hEKwHhx+lKT2ou1TiBLO5DRcAKCYOfpxw9pVjE1ABEgPL+kENzRdyNIRtxn8+T2FvfgYZyu8lPvO
4yllklkrrrH1xuF9Smifrjk/cPmFmXahQaP/daPRD+s94X+6YKYOPnVKLWoZE2gqudYH77PTbkCR
ekmQ0krxhUJudrsOSDo8TrbOAd+TW5jyS7TgsUUcS2lVu32B1m/ZlgntogO71JAR5j+lXvdmpu9W
tuNFh/NestL3xk2WVaqp2g/dn7/HaVewRU4JgYV89HTJj1BVWyt2kYyElDTkYBSEZve8nMw+i052
snKEh5IwvVzWDx1jer1xCFpwv5YqgwdoRJWXqSbnSInmgn2Se+GCqJeZL3YV8cAXPV+5ptbyxAjI
qt1ERwDu2BJ4xS403sVH94SmgGaA17x865eTg4XF8V9hqJkX9njkhsC/A8CD1TV/eSNPPlVEYf54
EQlcIeyeD4pZMFQXQPZG2rs93ZbK5DYehFOMC0ZMiBA6nJG4jnTiE1ofRQL9sqQLIMxEJVn4jCSx
VCDXJz2ypZa6jn65hF5JBgUjV/J6ye33zSQ9Uk3xo6NnXlM6+tukFqfppYzp6yTUFLxsUxrVXdT1
KQaXBytVvwLL44hsUZuu1kC0KlJV+tGTFXduc/f4iIo+GvJcF6YASMwAaqu8yet/NnoduyBtlxZ9
LFZGc6i1eGLIUCdjUwFbc2ivfihRIgA0lVi9AUHaQNxTyKGHQkRFJT+eMrLYQqzH5hK6YtWHUMd0
e2H3FuppaACH5CH/ZDc0qQfYNMRUBwPob/xzV+Mgm128vDhMWRFdnCmbMSNJL5JnhoVpcnyZim/k
cbTnZ/1188EY4/9I8f+qHATHINXXpB9GHtpLKR1GyrFcy5DB9etjDw2WfYZJ/sTORTK/o9kafoyK
kIyOvDORaRxZZIKGsRb2igCcqrPfSZMr8s6IFdEg7LzlDWJwCpuQFp5az+VHhwQIkxg+/noI98+1
4Rresl5iMfxxAa/szHQTNJy1jhsz0g0NUak0bOFMYa7kaRJU68b28UmkJokkENPY5Pgi+kwEqAbk
LcUK9pckOKsqYF6tMbP2sBi3VKyY26nD/nVI+/raObz9haXvZw5PLV2f4+/TaeHbXdHx3IglXlUb
CtDmyPTFvkEpr4WYpepe2ot69ogUvE/DRo879yf2XDIZGFnAtsOpo5WyHf8iDCuiUIJ8eLCtcQFk
A/3/oz/twmGVgx6biSc70wPK5pcVkvuhn/RIu19eF/ZbjDeKtVKxvfZckhNNqqykfsTy6v2uFc9b
k3rOrUiNTb4fa8OUXzCWwdfhhZ6aaARplJpCg2Ej8EUnSSURECqVwhwbwSU7dmkwHaVPnFs2yowv
ZpJ8wTBUe6dXUe3EQniYEqKoNg90nCgLswHje5MMNqCxK/KjzUGUSY7h/8GbHf4ctl0mlqbJL8IF
i+IbnilVTRnYcdvi47tQeIoVm9mnT5CNMFvxFt4QYmEbLZiQAeWFyuxseD0/Glbafgw4gzdUz8AD
q+6gOlOoG9zU42Da0fUbTtMnugC8EY6kduLfMDzB1ScbjqspCFYs6VvHlAwvQxKQHjZwSOCuNhgq
i5TOTR0f8KoPmjg+ImLpU8+K1hNefpRj9KGCVnCmwTV0JguBn/S4VdbP/8nA5/lA3fAUyq0DPhSY
dw6XbcASxOpAcve/idMUn0opG0wydwG2FRtfEYVTTCnTbPRL/NcNfcVDXrn8HSZq2mjWGrmRXo/d
+jtdb9HsZFSO1tCL2ThybXHYWZyFf4mfRUOn5gh7z1sitawlFnbjKVyjWSD1MHSj6Icm+mP6FuAL
B1MVA+4jcI8/j+apHl53rIAyvAVawf2HptH34YFnNkE+b2evHO2tCcAX+Ky4zD67vq6KG+27GAhs
6z7o9W2COjnNaD6xWUgbpiCUUgCKrPfx0SSde2rohgqf2kvbFsrenBTPf9U7uz6x2GpPDv6ZTPrN
gylDjIl7CS4YND3opWAe58LRQb7TCDh/ytdsZ6exmvkqw4dMqlkZ49xpAY5SqK55PAoJD3RD5ynv
Bo6lAFlakdOy4uXjkBkaKRM5A/KHrW4SG0PwbTjuYbmeXYgiDke8jaQZuGJWrRZmJgDSaXkSSwx0
uL5E4hITbJQLPBV+FXWsBNCesQFL5z4+hDv4UtLNu3CBa/4lJXt4lUGizCe7vAOU30ZCs8gwFmv9
Y0fOJTsBaDQUQFNYbxp2oM6BTq8QentCzyCzK7y1n7s3zaQLgQlYibdMFbJjLBpUq1P+C60JSRBW
h8G7UjZbi2gTMvCxCO9u2E0Jk8O9aECDO7rp15vWoWStL6QnogRq7wjxiOW7+c0dwHVJYhNs5q60
MLhKP2zFdGW4XPBue8ikKFpnrnnWD6eaWVK4KhDQevgw0OBW6CHCixY0E8c2vT4Xpmc6Q/ku7tM4
pzYeihG9t0dtC+rBjxCADhswtFxJq5RQdEjvyfr79lNjk5IL3CRqydKszQaIO2Qc/+qdmDBZn7MC
AeEvFZl6JIU7mN/cKCE5nCmVc8lJSdEAMdlZVv2VeS6D5J8QTG1xty7VaZ1CxqE8sbnokUa+yldz
jC02SYRMZxamdjy9UAiHgZJ5VM+5tUrO2dP6sgSfNa05GvlMA24KBkAhGJJF1uZXF92qKVRubLUc
kT+7zCAPFxVzn0MW9Wu/XfTVd8xTZ0xvte6I87JofnO7yAyRwyerpTw83YB26A8iWCgORB31bIZc
Xh0rBzGHxdfksG6stKWDOPn4FM6FW3/9nkQRPJjMDAavpr8YX8j9RKA3byVOjwhbNXE7ln+mVc2X
Y66fYPCppt7F59t3Hy2+WTSo95wje6sHOEm/8ISracBGyDd+bRvRMbrR2l8+/UuEbTYECMGqHOOM
dcNid//R/o0iVkuFOAKsTiLP9HGInp/Cg4vLawwWb9k5juoexMGCXQO15a2/SgpJNJfSErM2NTI3
78BMNrwqfwInS6vSaBPnwekGUdPAvFuXMBcAJuYk6KEHe3sxSz3pilc2CY2Uhl6Wofpit/mEkQ3J
JdUB/DIrk7IkG73FTpF5wc9/KRjZybxj34zOw90A2XD4PONrARfnjzEKXJADYudzZCVH8d2yr6V6
BGWINxRVtZrcP1HsBuDeNnIykErZ1CzFZuF6a8v8GMbgyvkWy7N0homi4mqZDieiDuFyzAjmFQRa
vG1VWBzuviLzazoGnL9HdLtnaUZ/dfE4iBHNHyx3RbBozbJ+04wnkarbXzm7TGwydFjDRBV9L/T5
fdAtXD9KPFY9/sbP9aQoBNBaWj0n1Sy+USdvzrIxmM7DBd8=
`pragma protect end_protected
