// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Z0A3Y9k17HCsCxObRcnzKSxNyddDGkjRrWF0e6PyP3PbEoTvmRKSXMe4Bz1K3Pa5p+5ihccBOF4L
V6UrbDOvLiG65qt1iH4qI0oylXx8HYUCIZ6aUKpzRJSbLk01rCL7j4HPEl9hQRsGWligr8ljKm0g
kQARt946RES1QxZAItWeLijhu4dx1h5goMLNOtV+PBZLhpZUJQIz9jHu4rWVmcwK8y+2BSJjA4U7
uTI4cwWzXDzL5fkBPDg4/QnJ65RXm5isnkcgi89cctPRBu/Xhoja0aaCW7ZZ0dtUrhOInWswktDt
FdIIaEWkwWEOfa0rV6kn/QNSBbr1ZQcEdgDm8g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 24816)
pgNF993C5Spe/FtX3IbHjVaqaijNNey13BdOu1pOTMYpDB9dOObqpg4hxHpEYDOYrTOi11zPkazk
0DdhCZ7giE/FQdMKhMzFJxlTvm52zKjrsxJiwPbYrySEr0t8POxAg7mQLcL5HxI9gAQgxevMVn1c
wxSQ4wU2F3ZM8KKjTlNLKhTFgGhW975xCYtewScqtcMkguAfQ2VnEeeLy4szKyASkO8RROdiO9KG
ltNqqK2V52YjmvXDxL5o1gdonq84r9VMJHADp+RoBJEbAxCODqEIgwbuvhldTgXSHJuXF80KDHhd
Sv/2aitpFeiHLnOVxAkaLWmGSzrHVMrFFaYbq2Ofxkj740yUDal+RnK9CFvJ/mJEMMrTGRt0yUa6
xGPRj1CXD036lZKFFsReDWiTdkM+zzVRYhD9EG2cAuh2CStnYk9SBlcByyHEj3IobJlWdargyYHL
Uue5SLGU8w6Td6ylNmjE6vLuvFDAENgveNL8JWq98vCZmEgUDDxhnCor6a63JNir2NKqQM3IDft5
KuqbfM0+HJf9MtXL6T0LAwyyMuR9kCgYNi2mt7UqwHAzQMJR9nsWljgglIraxNBm6hhHdNgJF2KT
YpSt3E5N6WCNbYaw3UWfx2MDZB07fx/cLaFb1WzPYnnvYXrkifcayeqzLsctmg2tjFg4Oc3icIZI
Jxdl4jahTpY+Nur220mW9+a/3Yc++Oajoj5y5islU17aU8/DC9UMoXvqoXUiSCRif9AdgzBH0aDc
9GI9g9FHBOAXdvSSARe4dFeELu9PN19w37odxajUa7VT6u9XAumd38fVqlcNUSxrfw4JBOyXuBe/
4Q7h3WbqDCL552+h50PmjQPJwqTV3Nsx2MYy0uLZXcMUenmRH/eZtJrKXXJ+dSp0+rIyI3GN6vdU
Kx0bE/GTBRP+9JgjZ7t899wDrEhXvBFg4rkmf3I6yI/P7NQ+9P9pzgKNLifRfVkH+58LZT95PeGm
5jNrB/LSd2Va4/LyY8Ef3Ic9vgkNwtg+43mnEd4Ghk0cHFpcFAjkRk+4Kx6Qx1bIrg4Ipqh1NC99
IqHudgyeNe3GcyOXCPb/cQk5ozmvMZlujUCABquxfr94aAvWA0gbClxjYMDvPmFAgIQu66RvE/vX
vxAr2eLux3vXfdfVA7/NTFL/CiPjeeEQG1oqinJ9k7afdCyJyCKThAuI2o7OElXPVVzOGEsiRG6T
3y2HsJjLonvL8h2JJ9/U/7dPBwRDjP1jwePAYtnxJJ39C5Y0TKSz/dyqIcEiVm9xfhDynMwQW2EN
uuCsczpvQ3fio8QcW9B/y+tRjZVdfrb5Wa9mjdJeRZrzJdt9S0oDr3bZ1eZ6KRag5UFWMBWUjhQQ
2fej6jQsY/D9epDAXVxkBv1wIv43HEd4Gq7dk62u3ZkAyEinTNpG1OUzuyiwAVGUq8e3TH5/0ehq
KBlZL6zlEunrTJe+mzDctR9PH8LXqKPYNYWXS7kOk7Pz46KVZvoaKoweqLIy5i+AJSis5LUgMXH/
q/yM15wFKcyctOV3pr2fa0AME1/ARcoLO7z04jiKtOOz0tbildlqXoFE9kds47ai/sB+0CFNWnG6
wkGvcBXCAMz0L/jJrGlDcHHFOKU2zcE9j/IvWkWtYXDeSpjcEzgX2JTsOMKPkK4Lplp+xpk67ztc
sdgQjrtE4VNLdXyXORVMPrrEaDZivdMUiwFRi0RDWXRH1r2sY2sTJRuROVVCINtkDJcXA+6UBlXk
sGPUDc5h4id6NqbpLqERS6FRlHXuW14Zp9KF5iX4r/9/olIFveqjaidotr8Y/F6BaXjYqaYhZbCB
ze4drto+OW4Ql6Yy9ZOTUZsp1Z2i7s8oAw+3djwUMftJWxddXNIGp9aUlOY2+NsFk6ic1Yws3eY4
DbBcBvPQavckfzEZ76TDk0S0yvU3+KlL847OJDlhu/16oiDy2mO4y9rvk61VYuGjcHgFncOzmN1D
QwpyvE1P45ZEz3gps5iZVXcV0i3cxL5CGVCWf21bmtSx/uxtbkQBibi1j/5RMQBwriC53Wiz3QUn
rMlQtnkjH6zujXINBKi/pp3WPMGZ5HQC2suDJiwRjf+5Q8rtUisP1Gn0N4H913Qb45a65i4Mkc3H
RsbRBdcEqtdaqEgFt3W+5XwSYQ1U3oIy/VtY2EoJuZH9WeA3ml3ThL0OQEW9vOtsQm1xXOsE+krh
5QPtZScaWQNBEukky/XJaByIAtoBH/jSiO5dGck4c2mkRIaGS91yGfrVHz2moo9nnEAfTtIemoaf
VhIs/xG0EfHiW/dxkpTWfXmOePDYfwIaOyjsKP2JQSFWLhwAlYFCZjgMMvMC9dv8zguleKn9mraO
DYsjGtImRtPc/xeJitDUN0g8T08bLOqyetIJ1C89gotyFb1unInYh0MsfWiYBQWsv9stM5joJfnL
YUQWc+v7JYeE1yahmunGbs37fIv9yQC56e5JpFFy+IeikLkBfkO5HCMCNmEfCxTM4wKciJVMIAXv
Q41JQkRYF0ZURN5gMdoJyxHeiK9EjOZ04FC8NrnlOMMZtuowlLjtZY3Re7frIA3mUf5YH/yxqsdX
qiWHgMz19m4aGjecf3R7p5Gfqwuw47Htyko6boIbN0nE0pkXAP92MJw0WQbOBy5GtZ76xKFT4gwZ
BfUr7gpQOezjkBpK1+cNIqJ6+FcFxMyu4aMv+Jv1S2xdMN/tCXyQ1AW5jmC0Nka16B6tFuRhihuL
hlYAZ7r9/A2BAVd+ZaGQE9KvUFr//9oCX8afxTLOAYLApArINvx6tJz7YOMCSqRAl79kyDCrnLpU
kuqSU6UJoKpttIsaub08gI34FCPe2m9ynBNnJMQTLpIPUd45OrFfUNQSSQIpGkToT4tQAkOKDBpy
2pVFtWsz6BRvs2mBOPMVFJPW74UN9X16R67JAPt80iQnuDj7dwD4sTX/vqCpbrOb4KSeYWaASF5u
aETQQDJpLDlvHMfBF7647N5jroMBkFSPIfmB+y2BezkMkoVRj1eE8bpmbhW6JiLeMg36XXnpwN3+
RQzqr/SiQmUxjiFN5LALqwy5JUGh7vK67SglVQLixzKCBlMsQ6qyoM1TR8ufxQ0+FZCQPn3c58oF
QA0M33np/j3vefXLlgRoCQjKKvLhiTORzEfRnZFPcXSE+eTmQPIe9DWLH9LuDxOJPWTRzAKBe2I+
ZkG4uwMDons3UR3QY7It8w/NTWczk3gZZcUckUzL/68VQ1xkmTE+/D087QRimCCa5ZinI0HKTPOm
F30BrhrLDRYY7KgiEaMQYg6d3lp/9dqPoUj3+tdFnY8I35NmUMqJalE4u4vQ+via5TYEi5PvBYz0
IBZA/Ya/sP4R7pkwpsvlUuGygoU0kr3CWqCVxaF/lTcLG5DFYqDdz/wnITL0v+pIvtTKxQBk+WkL
PvpVtnqaRNa1fakZpdB9eMahJ8p9Sj/1mWIwJzSJrllAAIb+6QqoruOFAo7g0iJ9Y8J5d8vQnpZ3
XaApsZZdTffuD8Ko06xoJJ/ciC8/qDCjcnOzY6pNuoocNSVJCxKTZd20z8A8a//1KtzRah+LxaER
zdP6GD6pa458WzY+hXcBurXxneaE/tR8BhIefH2xg4ZXCwDhjW1O5idsg9XMuh3RjoNq7Kwmp1JI
c/ZwnQhmJ97xjtfuTVmOGSrnxhxUGgiQgtYd8RFTjdnbAhot62fJuGfqdl77rpszAre7O5zSndav
Ifnc5KUo6eAhN5LPllTvIb5e9KH8w25E3eIzPxmnhEUNBsyLPk06QBQayN8UfId5BZfs1/QJ/dvY
shewuuqUPN/jFqdMJRtRXqQJwPDPUApvmS+c+q9V2K/z64i/BtLR10hZ994xCKINt2i7bFBxO/Ja
vibQ3z7RMQWFOcdJsO8o8tw4AAO7B3L7F9L79+MjUUTTJwHiDp1qUL8363sZQYTVEGZVSRIYwDy+
e4M8Jrdl7Cf8RX3+tmb7ZXCsqLe4KuDWwDIPvUDh4tOkW3pxPpCbeCLemNYf9JcAnM10w7bU2/yE
rNIlZf3hCm4k9xQ7MALEymsvXs+/4zForU9c81jQYEn6wRleVG3kv8Wdgt4j1e55vAPj+4thNLRh
Vl6/pN78maS9ILT6p0jW7JduLwKieP1kJZBoMck2TXsP+mxyGc9NyrOeJOj9wIPirgc1lgVquop3
XDQKsQvBFsfbGqZwjB7j85c/hEdZMlPc8Cn0BH8VDGnEMU+fqUUSA5d25blnNHhl6rj/VVulJZ5K
AnPEE4RzZJOiTIP0nrFtu7V5l2PJxrHEblgubXEsnRg9PokMaIICs3s/1qXWFK8Gx2w89N0wXkmn
R1vvVaZPhmfyFhxKac5bTGkiS/gz1qvtLhudIsQl/1imlF0o77ISAFptrtTChJHSLscDWsf4875l
YURf/QdYOkv9M5mOp3zcV7WpUwG8z8HTZ5cj8oXfYGIXjDwtiy+2kRna0f8sgLy3zlo8Klk91X/L
X8PP9dtCv8E4l4PvJAIXnttwG3h+ookK4s+12v8A6PZCL3OywR5kJ3oRnQ+IlzT41AiKArZNoolJ
6gIws2rW1b3fSYpp72NfyziPkZrABVgmRTHBbsfmKfR/+RhuKdnoQfXQx1oCM53l05u0H+9Y8XKf
/GdNlOgD9hnweW2AhmQlCiZS3/LSQHFIGdJv4vRt/2TrC5gifCMCo/crYwkiA7SRmnmCpjz5IggX
IgM9CKn3t8K3tgTX36v+vi5oxwgvY1HL+Z01XqqukWc5r/iMJp9IYym8ZI4T8doT1GrUDFVx+/8V
tBiReu+ifCZmDW3ThGAB9Kdl1kKYXanjphn4yHN3MlSfen9HUqYvk+t0cpUWc4GwCtSZOj8/OShj
bBHDWN4/Xhrzpxh9ZIS7e+Ovjw5XESF00zFEumkNzpOozL+TL0MS6Py5lkZzzv+WmhgSM0Md9zet
MlSV06IutlYrG4F4DK3ZDNmtBxv62UNm5Qg2wzX9nI51wPiE+mx1oV1gnwLH1jaSuvp7MGiUWWNr
FIIOwPPnFbizJkfvIJh+Y6hkuzCmXaYZ7wjHmSfVFKRW1wjExrV/p+8V2m2L2TpneXDKi6m6HmLd
Qpg/QaQKBLhqVOBwIgRYt97ku/5pY7g04FnWQbHlmM0egAz4uMDSgbXrfE8zOv1gO17z1yvz2Bm6
luNF6717yaARI7TBEpc+OOMns4VYDvIBMxD+Lc4nDGHr5hVCXa/Qe2qrfMUHO5BYHGjuV4MtoEdx
D+7UGeGGLxmZ6JXX6PV76HqAw3jVCIJ2wEeM/BsfSlDn3g8h+3IbLc6vHU2r6JU1nfovvoxfCbYS
k3MNA/Tih4kqX27ih62XyWtpipKlwwr79vHDlcsTVbCUCttNo8KF3toM98k/YWGy8BowZTz05Svr
l5u9nzZO96f6CD/wpULhVJVx6xYIUoOLV6iUbA2mGRPu5iMCSM3YXjP+6Y5CvBkDwWCze5X4tA97
d0rSOnQdwrrxMx8Eo22H9iBY9/pkKYZdmhFiHpTNuOy7liT30nmgM2bZjgX4WUtKYpyaQhsy1Qjl
Y3YHdIUtcXGWHQCXO83yySXiEKHly1UCuX4NYREKsBjJ3M31+Y2N8LnJLQMbNjUsPAK9xWUsDzMD
vw2muZPnMTl5NwgTyl+lr5l08neUmXR0+VVSDNFmUsOPlhubgjub4HMbEvHo64s7S3VeJpmUFN/h
cH45wmDRf4/DxgE2wKOpO1Stn2EuMsU0NTFO4XTYvtOxlZ1VHsRqdEAfqwJTHH65ij/IZ1PfDT56
2r4HIZo8LAHkY+IN69pMkXOeHN3POM7pnVsHMoVce6HLApLzD9TdWzL6wd7s4GzuLLTxF0jnxqIt
XSn3lVqm+Mf6imQxQwT683pJXR94j0XrkuWn1hfnADbPQ0wSAmyUIQ4mnagtagzYtMhw8fwzR5lT
rcpn6g1MRwcsCq1rPC2pSEnTvN2lZgqPbsmt5UaveoPkch82PVDGig2d18Lk0o2ZMaPkn7i8stva
uY8V9EThzrWIlGu2hR25q2E9AzFUO8ZF/c6BdgSUYRKdSdeIsyfN74BvicYfPe+7VA7UtoojjGoH
XJAtXGqscGfJZOhZ86zzW5Vz8GmCzrhtNezit2urO9dzWKPa58l3FYi9SxdLcSeqSvpgl9M61kwW
iJZc0LjE/O/tIO7oRWBdegpiCEuNxYoyrDwkrB/1hHGZJP50qYQgqp3994RgUOf5k8+TzoyMmkfR
N1qXYRsUGVyNdkwfP6WGQckL/ft8UxE2ik5ASAOS7TMZTZZHM4r6RD+MFqc0fd87uEc9XGWP3m50
KOiAYxEvcqIIMhGWfHydIE0isLdjLZjZeTVAAclUN2q0w1oc/12QPsz/c319ANrpVy9Y5yYe6edd
8Uk69alwD2gmTZATlPB8pOcdc6vnlzhjEzo3s6X/tdisT87n2yKDXe9c/8D2BDAOWz/FKE6AW2Se
fqKLJOBZmWUeRMYAurufgS2qYesCIzVi311U1x9DonpR7JX2ovUvBVx4cfckU/hvG6jtAFIDhitd
4QW6WbTs6mFB3IG3M8vc6Gf9sf5g7ZYZB9FLubQK4PuuYAj4MkGPP7+SymjGjVP2CmSzrJSi9rtm
jNKMOu/GPDn/7pTCC0M7B6xK9PnheQbUYAW97A7lnOaw4pnxkS6HMqPLjVNFApR8p7B1XJIQDcoU
rMgLmBsn8us6XEbVZj4XdwmpP133cewP6bG1ThvEgMVpmtC0K64kzP/9iBsaxxaqBF92MKlOa2r5
Psb5AxicXmE/p+3xCR1RcfAb7kiHvKbg/ZUeoRQfsmZJKGjC7Zu6Ji5o89eDbdgdr+GMal+U8wLK
ZCmFBLedNi2rP112tjEZ06iXCurY+s1hQ9fTV1WtarXrt+kBVCzIQG9aumegk2SPxVq4fAXGgfcq
tPApkWJNsBjS9AI5npzb0RAlor+OdT21ZCLea/W56L0L7keNZxNJfhk5yVohQRaGnIx9js7zgM6q
mxqhiUWMr+gFkywp72YR1Oyawp5w4YwZdQrN1x9YM2lmEd1pi384pGWe6cjtSmeNA+lIjVar9+SP
BpXOs333oP3Boi5nuYWACyp2NRrwmHDhIssrS+ACL39EQUAvLmEjIHdCybk+Zg/PXEFg2m5LShOi
Cl9waEAsJ7gAgI6sP/JjwTc2qyM4AdgCPh2tP9mgwoSI8qjZzBmVE/5OZpcAndTwU+Z/XknaqUOf
BffIs0E2lfIjROBtU9kzMPVU23g+Lngwo1H2ejI+x3c22KUyT1sFo4xfq8kVMvbmg0aGRHKInhCQ
DWWb6lITMFPaIb3PqInjRsxFiIg6ttN+nr2Qu9oaLheqCcTOHB0gp4Gpc1teJBQA58G2GnnLIAc0
9821KhAGVAFcrOG/TseuwiA9dQTQojxVsl82f6RNYuiH1ua3jIXsvL/9g2QXOU/1tETAVOuYb1mn
9V1rEmcu3i0XtdzZH2uywtPComTny+85iMWaV17JytQ9ADB07yPnZwitilQ29lk6QSCDrFem2NM3
78Q2rKm2z3zneCti3V2CDdWdkHB5a2oj6xi5FNu8mcynEZSZw5Pd3tlMuCDnzY3DyILItfck2Jnd
UkLHSZ8JcFEY2W1hMVXnml65Bdo3ayzEBwphkYLym/XUUqEZOCf+7Y38Aq5zVuIK4RHo3Xy9YmZr
O+VCFVDicR9RGrjCBV833rtJ8aiN5tW+o8PU81u/KEmdaWc9Ate2zJL5yvMgD+YZp/U2OA3hHkwq
Iy8cy+Am8s/JR2NPWsR5GG6qhtFVWTomU6Znr7bVs8xg++N9NhCqD0EBiw9C429Hg5EHymKNZlNs
LthmRHHEzFjM+4ypubvukZs+oNdMjuMPRg/x1TgLUgcjLhZHLbLApqQs2nkeEyY2JsZHUAXMVmum
y4/tFvUH3UA2dFqrEZUBrxaEiChnOyvIL/nSDj71xmlbPpD46t5t4ZLLRhyLAUIKrXD4uAGQGVJP
6tDWqkDAOYuD0k1pZe7BGJ77Y3RVGtYvFjEgEPH4LtmvIsVZiu1luRCBaO59l1QiyNHfVhMYtR7A
SYw1YGwEmr7w+go3/wQeAV28LsLqe3LVcOIp8LRXU/Rcajg6juDVI89h7HEfP71B4CpOY5lA+KsS
KB8b/6Js2rAkiKqDUEbzHkvJov/gxQe/mtyLxGtjkkDZ3MTJ8uib71rZE2K3136mLi7L4angiQ2V
Lx0XX9qaKHBVGU5oksDeayfSGFMkw2HsExIzHVUWxJe+ymAhXtMMgmwyW1bufxQv6w+o4NDSl05r
9rK46HlH9LdKMfsJXJk+d5w9y3aHPcr2lJnhNFcY47gOHWwiol+1ZDCoRo4mNkxzjMBXtHTDVHDP
NmwIyfvV11u/tBpAbMaz1W2im42xRmC74aA5hj+ZGoDIbt0SNBgQWs/kQoVkr3rWfzxFdplQjN+d
bMx3INDcU40bjwzmZFcuYGl1cbaqNhJA1cScz9oQnc5NdTOCDtXuhBmOSC5xlvAy8Sl4OUNdbchp
Vt/XYC30jSh1CTR1Oo9aPREDNkLdGAg7F2JhYv0JhnFZ0lcVznOYsDzRJxUt+t6nafrafky5pUxa
fhiJ1TWdzcuGJOfe9qekroYoWJqzKNoI+yxmFfzRKPhU4pzd3haTODJeTrgUo5Fn6IO+0FHid2kE
IcNE2K0AERC/loy5eO5VVM5p9lISYz0plJ5owEGlWEiUETK3H6afHdYYlTfWZ4ROh4PGsEr17qAo
88Kp9jhd57DK6amCBeKOxGnbAHgidtZA4DKmsagl7M6QXAZfM3LkhT4+th9XT7y1++J5Cxr+O+OI
SWbO9LK8R5Q3hrDXjeDUNhx2Vz5XW78kPqmXy2Up7uHCv/g4GtInha4o1+gl/YSsuOboxynXcl9k
TP9yE8+WdwYrjOtlR7DtXVE8Zn+kyeAFwaQKwR1lgfDoY4Ax7utEPbpdidKdjL6008YDDhcntwXV
4/qvoqFMKFa/g0HM7fI/xJT+bHT3tmhpSYbJZAq66NBo3KreCSt/Xx/B3Gc4RAEHUB49uLPGKD2r
PHD/EBv9N7GlzVgWzbZQs5SJ8Aknc1Unc0C3oqVKVjF5qUnKfSW5VJST16ojrP1HfzB4g1DM70O+
0f1UiKtKhTVKPVjoCq/JMm5OkCVh72igpHlP+n/Ku0Wwpy64fZsLoRpaysrYgfNORlkbZhD08Tk8
H/rTLpdGm6eV442a7MngCvDCNrroXL5/G+RLRqXD2ANI8CUIgoSqPLhIqH+kuen1wAHClxBKPUmH
8DsnfdDUVJsBT5QKlfhWr29d4pOS+s3EloXF61JQUO1xK9BcFr7UjL85c3vExUFFt3O6qLXpJPPD
ZDLbDbnOy4zQj7RmunF5BKoEeT3qCx63nRytvNVjKNup/3pgAAaFO5rdbSSZb+aDAWQw8dhU+LVo
LBF80Y0PHTc/vS0aLSYqXuFLUmhhYTnmMxoCzbKGW4prvUXY6KJtWoaJoxpUunYgPNqd2dYU9s98
NuyQkRG9Zu1wU1R6Fufbpb/0jA7qkx5McqJbTiYgdolxoBwpoODIMl+ZZnhC6hSEaJj1dh1zo3cv
Q8JWngQ4Jn/0Q4JkyWgqK9h3Ge7bZyIC13HlSAJkyfSgIdeOhESE2USK3y0hFZTjJRAW1wWYP3AI
6GmpMF6h8qsojk1vY8Wntv11CWu3wMMES0+5fgtBmgSrPLVkNFolrQ/m8nsYkjaIByoHCi6vpHDv
zjSfkdgl4MdLdwXKT7lpgKkYoPE1Kn9WGOtFHEzc+YDCnCgli4bwvA85fIjt/O125RflqwGQStSK
WVk2JadQyVZRnmuF98ryF7isrkywaR5EZrdcHKYi4HKgM2mfTga5IY+CmJiOHSabpnkDwzeUw6/K
qo81mesQezQeHQRps3VjiOA0k5kqZa539zhA5HixuMA8Pv3VD5AQaWTPz0Utg4n8IMaI0ng2VbbM
maT2sSRR8D1jhaI6toV3tccsq4KRQUr3hulUxFs2gE1DVpguxsWh3y1rLLsgWn93f9v6VMtWJkkU
05Gpe3mHpA80h/7mZZX4aut2vWlnZu1ss5X5QpGNFnz37MAqgpeCQHLNCfkjjibUlnyDO70hC64h
wLEJrNBQRQ3Wv+mvCxTM3Fn/qUDS8ZWf11h/ZAQy2ik5zERHKtUQ9AUpVqdMOevPTkPt4v4Ffvh8
LwpX4MEMJ32AQ32SahM9ht71ImVrfU5ZMwT+naKrCPepUxUn73kF2RuASU3pldO1xoKQkHPX0stW
U1Qc23uATKa0WMnt6191MMk0KR76P9SzMqF1ITMY3i4JgmtszcroIOufE9S9sb1gizc4YMqMl8g3
J5L6MTOJH96hiPjtPUfrtpuUWuppHp4tnfmfjLD9ISwsem3d9Q5vkWQsPgYCXhvXmU3olAlP+E/G
pN/V47n9CMzTh8uxQuFfrTRgECb2AwqSvlw6eUSxb+jXeeRRGQMaAnkeZjO3Cujx9+WYTe8qjzS+
REc9Ch8oBmYwcddt41Zi20pm9nViW1lXt+bgXFK6ygDMHOdNuvJbwNIwBudKXKtIr6rKRxN1S4xC
+M7QcNpVHEsndzEhtxXcEbB4B4Ji8CgDUEzImxu494cvAx87sp+AqPb5TgMtjaQ2oq7jaX1tRvNo
jXuP6c+YX9tQR5rzi4arG4GWiivOBv6cXKcAvXsEuvTV8r7wft8TcXyKh/5qHzTJozyNUjUUthi3
AUfKNDlCKQZJlLlt0m/kx98zZG4TAQL90cs+KEwToZfieDPrFjRmsIYgfYAlXZm0X7fnHr19rJoS
ABxd9JO4DAc5szHsZEsKR8XWdsCIPYxj1xD7iTDwgDRVSP8nFFvuCqocc6i8Ql+wS1Hk1SYs5wDQ
9PdJYxHTD/hTCxI2nGTY5r9wW0ZEIIaSsT3y34suy9sJg0BI/AZcMhL1M2ZuFQD3iLI4mFsS89Hy
qelbHIvUKQjtv+7GjGQPxb5Hrq3OlWzsLLWU6bvGyCq53gSBT8A5v6yjAS8Zq/1vZ+oDggw1VOP4
bDQ+bYrxyzFkRGsmheM6VV8tBKwVzcYwcXVQr4CpjbeFwYpT325Slmeg0Lwe6KAdzVMJMuwHxtQn
DqJLx4gb5UEgTicNmnYhwn8MbyR0unqCTnRgdKM8N1R701o2ho1GUeiOARWCrzdzk0zRq44VgPZD
yVPqjbsAhmkfoJrn6zqin/2hnQAK+nHoR1N/1hExBVpbLrsjjGkt4XtgYJJD8Kfa2mUhHOfVJ5fU
UmUllHm7wQNjkwAZX+yg/zptI9x7WRU5SbnC5DVTRhnkDFYyXQ0YLNkBceI07Q8tcaa2yEI1/9hi
+mZeiGqX4YbwXjzJg5szNzGwuvdpXBx2jN1aRsxg6XA0NSWdUv/oa6pTplhZXziYdieK/XlcxiBI
CjQk2pUg0SPeWr6FH5Aeeno1Ny1ES0FIf8j0bA/qQWf013w0mOUqf+mKbXpH2N+v8Kk9K0aLfdhF
ALFJYB2vn1qKwLwriV1JQ3LnjyRqRLTW+L/aDfGFnEb/wvPIzchzYyOl1I4mAZL1j/IaMFs4MeOs
+qyAFrR3yoNiy8J53wqRgdFJTUb6TWFGfeGrds37WDQXHgGK8wyI5rts9oMFNNxqyrLwBh+AVqMJ
I6PXKeLKWL2DPKmDjviMS8IneHSsC6SKPaHTi9WpnkVWn4QrRmerAJTjM8qGUWPFLkijdIV0DnJa
4rejove/POc4wDBgJZzYMNuVlpamQG2Rs8eLAGEEAciK8+UznRPWgR8SghCkHYsLiYud11na4E+w
Yraeb33yvfLv5cfRtQ6rvwC6JECEG3biyLiv6/tIfHvqUJnfUp7jZUmKmGHWyCNo68qYKqClaEpl
okuSD3CTMd8R7hb1vN/F2VZGpr+OVOL68PjrNSva46JsI7daG7u2sLLnypiwAY5kFvL7oM+jW+q7
nA77zt2fepiJQX0i13hfmbWDFCys4e9jFpjPwRairOk9K0U+xn/tvkbAZJvtr2nprfkkMdXEPaq7
CYAQpBpQTfXNKzyrsqi6o5VQEcFwCcdxzVr5PvYizcwvPw0Hd+jSRLhV9li73bf1OgE0qSErynpp
LYoFrALouTDznPdNRvuYMAqJwhXRYmKJG9dLr+61LkkYVBX9Pqq6tdFWQHdMDQ/KTgzL8AA2hKuA
lh6lJOSDlcDbhx3KioKyIqKeH/JwRP+WsnKx+MvoRBT08G3nczp77TJ2rthwRjc7PLQJgwEMZxH3
h/b6pCvEnNYvvArxpQeAVzBzaAQGVqdAX7+1zgoZ5NNS2/HP7Fn48hzV/8tzN9nqDLiGtEp1lkBT
JXrgX65AiuF6ji9vcYtZ2Wr31Flcq8O+E5tkOoUGB6PXmwv0BA9TVYqhKoPz+k+UFCeXb02nHV7X
hLCTrKc+hhwi363sGnJUar602daI5gsbZOClhtfG7CoJsbwYJ9mkiOkgkjSmEzOB+95ekvNTSMdD
TLlTCg/NuFExkn7aeA9SisHG1ZwTG2cZDiM/9sCgMMoTn5mlxWlu0ynTsOTVnhAFjszHmc5+y8n8
p3FQALF1zqZPDNDFRYW5u3t4bu8LpfVrwdv+EasV32bG9Iup9R703MPpIRG1zQdJvHf0z65ETTTS
ngMIhb/9DvvExSDK+i+lxGJ6MjE6ASxooYkUGUSVLtfNm5JeBQzQdHSdlwOsoNRG/bDXn2v49ote
/rGPLJtRZanwHydYFSTaDX3u2PP61HXksLyAICCUL86TSSdsXeU74vzTxVLY3OxWpnifAFDewDoM
VBxuXP2nahejM3Nd19QePfMtnChI323P6LL/fzQKXwz2+gfr83DF3BABuOz+Cz7LYNmC2j5T2cjS
puDrFulBt3i8AUG7dbL+wqpoc2SKBt2d8arLSGfAL8lER++MQmNtYNZ+ckusy+z7W2KLJ/hJA0Fb
rBiZaFYRG4wvsJcRa+1xvCiiys7eHo2Z99Q9HWe2PiaOt/ztGN/vjUuNLin0jcz2JX4OgqS+wyEN
DTNAg0XLn5DvCcJ08uYknai6FgJVkM1BtbiYt4swA+in/u6u8YmOAfI08blPOwVTqXrgnXXfTEIU
hFAB3tPpEYmhLb9uBOVXF2UnEF+UQExKqPBKhgPlG5DUR0CowElfdF19IO5o01nyySYMXay67T2a
jR3NAV5W+YcIAGQX0ZT61yrUlxxOXcSwEanpS9e0gntMB/TbyvRk9Ilm5sCUrjU85EyegV4gbf9I
4u/V0W1Up1mqnj66ayIMLU0fZLQgl+jpxsVYGbCUCpknvHO1uy6YFkndERIb/CEcAgDn279QcBzd
jR2O36mvN2LSypcef0aSR+6ZzOmkKTPMR1AUz1RWwA2s90WV7bSFOkwqrBCMpvKBUQ+m0VtG9DnA
U0RNvj2Y3nolAsoh7Ab1OFe9EF90TNx5m/gXWF4pUb792TiXNLVg5pJJvEzbMmJj87OKgvxz2V3R
mvouGk87sluYjkyHjGN6GSSyq7PjW6wUPkF/6VuWMSiJP6aXp3poyhYRWOlhijN+K28h4IzbkOLl
zi8Vr4AcM7JoHLWdz8iKJk5+ItMxN+afQRdrFfxisTpOKCriwNte73lTzRyWLp1FqBkYVskVD6hL
bU62fZsgrpA5HOaP36WTN7gRL32Zic2h/8km4+T0Kxq3mUb0dsjprJkkq/OaqfumoU12HzRlXCpX
/DdXpvXTrCcAhL6huT+b1WfFpEqGRKLPt31YN2vbHmtqlYCK9oMw1kDYiMbLCgfuZyW+fJRXMix5
O4yxakFxI13dAh6DYfkjqGkwMcan9QWgNW0KWEd/NLQ4cEGINDZiAeysk4BgjX+bHFoGXVD05qNS
dNPqo5LOD/RR64qh+oHl8BjKLClCEbmXw090NRCq9MCXO2dHvvuJAh7SR8eGSrnq4CTCc3oo0qtu
g7tiqTm6NWiMYftlFx6phThGlxp08p9r+YMaoWYPqcGE5z07kdyqhTHYg2c98x94O9dxZano2TG3
4qy05qjjMcrgi14HuOnMKgt/58UfU9fPuphmRlGU/7FGojNQidbWkcWfuu/LCh9d1mG/dlOQXkna
ahOAk6KhgnzOUXmn2orn6aB6hdmwM/hkg5aDUvCoGndPc2N7kUD2h2DahnQRaTRNoR+6OJk1rFXu
wHiRCrAvBtrYrpwH9ueFim6VOAl/8Amie6oX1nCKg4rrwLelQJ47RYVWcv9hFCSn6ERVK/P9jibM
92WWbAj/DOA8S34cgi92+l9ljdzwcUsQoD26YeEyqNL6sBo5WQV+SELgWdVGOcvJ9jI2zNGtg/L4
1VYo3iL+CnyIYlZVW52sYIpUYM+SHN+pWHb/4HldVsTKZh1Sub/IK3WCulQ1xQ/GGtI+2xz6/DHt
b4CIl2TDPKzUDxbsIBjpCVJsmrCGe5HX+JePipFDqDJ2pIgigEXk6NeUGypjpeyRndiuRJ1sluyG
etsX0m4BFfRu4LwebSLIjBFuPVXYSsQfHvypd6Zo+yGycoZkJSiGyVom0pO+U1wrpYKWIOXYHQG4
L27aLD+6xJcv7Z5lLK60Z0+5340X0WdZHA+alb+8DQ4VtH9j7TPzSibLfHIrWxiqzWqCscgMOvMz
x8muQZVfxoJuJob5lzTTdDA56OcpmTZJL3U65xF+z+eZu9Ob2fqMRtHDLP6Zk7OY8clF7QWFzsn/
rFgew1Iso+lUrlLJj9TEkrK18bPTIghMF6DlavtVvzOHfnRuzWcSmyHdDgkhdr9qBpSz4RqVNzgm
a7YiIXlQrTO1HQLzCP/5NzpTlfbvuzfHxSE8I7o119AAgpkfAhDXSaXO+T2XFY/pB8SxBnlxQjYw
XQw1XY/1jGtxE/uG4Pzr59HyTDYV1iCI6Ae0TzWLw0Yl70M+jiN5lt3KmeV/cVIMBmNO8sKPfhqV
xS1IHk0jHsgreQVb34nqxHz37vWyJr3WOsx/EO8nEI9kMHSj4H0QzvOrTaPxr5k5mvLX23WSOLsb
SFBw54YRexoGBIT30EjbFiX8KG9No04cdtPPq+6S96JCMA/TBqUjAV5qWm4CbWm5wK++KDCuyk1j
NiG0nGHG6r/zilq6ZiqUg7Qstx9/I7L53qjNVpefUeb/iYNmVfCEAl1p6dkdJXX/rdWobEeEVkkH
suGE8ToWCm7ukDvT8AXMUqo3sokmbKMgjbBPcoPjmEI98sC96CPgn5MfZykLAfl6fkbk12tAFEMF
GlSJXSyyfLjV3ZHbqfXfDrZFR8DO8mJtRUeQ7ZGDRq+O8kRmHpBtB3jWL0+nMZpDY4uPjQYDRtX5
Lf2lEji2/RT/jjHdNcc4RlRKxkGblAFMFcwEZgDuwxgo+LNdAwjEiDJFm9CjXEUW7YSYUKPQVPvk
AqbdplhbAZOk3kOjDRFviuXxE/95I34nJTZAljlbF4IUpLIAgNO4DXMW2jg9+kYAjDF5kEtO/07f
7yisr06ogzLXGMOmcXtb3y/fSxgP54TqiNZ+weHJM6TEjwppR9u2beKbo/yleymXqAMeIoj+mVs2
hM65IK5zGHuDTmbjw6WgQkVJ2UV7eROPf/tV3UtA56cQLc6HK7td1jbkzOKLGKo0aS6wkjpRYE3/
r5TrNjAdMuxqxsscvCS1boAO4IZHF7aTXmgn/1Yw/tX8ThahAK4Yo2QdmLw7ePE5FyafhL8Ga4as
JV1T+hGd56VcnAJDyjiRiK6paHaCSzU3vGVFk36RoiAisEUngP7T2iNO2MTrM9dwRRzE5C4f/Zq4
YcmqJ10Pgt16cgCJC455dxOkYYopRV8CpJK2CfqpIyApGq6WM7C5FniT0T90NwM5jHS8df6puuNN
ZnBh5TpL5EzxKxVG7bynrvdzQxXOx/wPbu8qocrpUUkzt0T4zeq44G3Uy4gqT9PPMFPDG9PwwwbO
RFTQrmMNW/yNxH+WcgbfR1tTTNPdGwxCAxtmEAFJCORGp21dt7Tany8wR+CouWUWc+d/pqK632m6
+MmI9J8dw0pytR8w/EtvhPvjFGrg+0zQMpBt/85quGKS+6yM1gfhtqERDOhh1kEfHx6g3e6VEUY6
Hp7ZKOq1/GqCXZR8gLTbxJzDwlCtYu9oMx9f2bD79OcnBfYCI/b1UKCZEO7XkQVD3z+wr0TSq0E0
yvybuPUlTNUo829Cg8eWO/BK+HGTKZnajCHKEfIYf1iBBu1/jTraKwZufcCk6d+VuGVrrgMgDkt2
9jP7fnl2wDzn0ierADzV3gMzKGfe8kfflqMQTI2t/1NLMn5wadFDX0EDSBrCh5x8uwNYWm2Wmkq3
zjkbkfJTtXUsyffaj3RGumT8x6PpbevogZIUGvS4TzQSQWd4lUDsXfsyPGCUgVYdx7S3tAbwz/0B
HpH/I4rH+qqL3o/nJ/v3PiKxf7GtOwmIFfQ1df0mhZRg1ZczJzW2vf/ItBlIu9K8lDwa9WyYDu8E
xURCbZFAZi9SL4EYE+ITjaZ5i9TCvMWLezYOBHAlASg5KpXrxt/NSaLmu//4z09HM0hgcfKWeYoJ
CzDGOMg5kdXecjKbUmy2J2bo9FUJNaQMNp54dzHBXi4EcUouoTJZ/13N83McbQJWw8JCSGzl5hnJ
zhnqZL7ExL0AVpbUad7wAmpA9vn1cx5xW7jsrrLnqIowSyS9dMUemB35Yril/EXEakWgWE2DjZai
bC2hL6OO2SvnDBw9zAVAgP+PHMpR7XtPVW1lUWi2aR1bp90R+sEMnuaUfbiLNnFZxdLsi9l5XYAd
2QXrMxJAMhsnIr4kLBLaYgA2YUWgTpruZvTWIFQxo/dNenTM6a5AXHtdIba5UzHpWukgm7eN9EIu
Pa5xEA1j5oQkzgObWXf8es6lXoDe3dNZJd6RORC18FlQLimGeD3qCTyja6SnrawMDmNR+f8AsgZ2
f3zkvhNYbBE5qDcXkeI9LCY5f4MSNNAPbLpHlK+3sFbMcIbWbRIRWT49G5wdMp/jS74HyMSv3BGB
kgkfuswD4j+UPgILkECamNXsis3LanjD6cIU7izX8FvyXDMncXbb+P1yKTF9OF9+HCfNFzghK44d
4yaQMiJTgI9hYMni6SsEgV+WxOtWJg2oHq+d0oa1ejLdhYRWGWqCqByZuukYlji4Xg06K3gV5DZA
d+zum9Df8KImV9P7lLw4uLJpF4aNxWl3nwsSrlGbpmtcF0ns87iMrVX603rU1/8EchodB0B4kswc
hKb4sZu6uHB0RbdKep3Rc2S66YkmM/LopFKIH42N/V31hgyorSAhUwg4YPM2sqxKO0BvAUArFlt4
Pa4LPhr6A6e6OPDTFBXnzUraxQn2kR1YFZHhUDDGQfXOwgkaiE0jSYWqq5o8CYeWPulkGk1oYgrJ
VgSYpl4UhI/dOGLDVb6xDz3qCzTK4aQcLJVt6HVzCC/DS1ucrqqb14CFxIjGQt0t1q/o8etCrnVq
eW2rsDAsBCoEzhH5vyKQ/7dWgqZC56BixSW8V+GxCVDXT4rnZlEu3/cKFr8Opzr5ZJx1PYgUoC7o
0HaK+mZEGmim3Vh3EW7bFAJbA7w5jZGyZ8RS6GL7HJd1KkWUzIg/YgKzPxwSNIA3kAdtcmNT6RFw
yMljA/MhJuxGQgIU8wAdpqgmHgQQQLFnKzhQIUsad3A5rtaS2IJCOwJgofAAZNKhRUzPg6aOyIpX
jYb54wsrujMQ/ehuYhjYcJxQ/vWRhguQqhJPUOxZnpMgLN6fkU5zzfBgTw+Vdcqg5OmCSbbOJkCb
PuMBx/RgCDCOwP303XsESZnlihwKw16KdHnCkZkWdf4zEuVyXKmmhCPWrRUJETzxSaGG0g8iWL1I
y61Vl8+8rAhpmd3dbo4HqIZCsbtbz6Xk2TvX6Vs3TTgyjdsnkXl/qE0FrmYCJlaxB+jnGtasaQ8h
fGRL0lswVPEeel4qGqQK8Ai5oHUkdekTyAIaOvghRNjgz0OeHvGlBsFTXlhtyJ1WYXUzkPdteJws
rJUk1PNMNR45fZOXdcbH2IJynraNElTP4xlun2c02OdNaTa3ke+BxJyIhoG7ZHmDF8RmH+GlqX3S
aaNOIgyTwkOopHJF+vpW7WGVUuCmm2+1eCTnLaC4EsqlhNW5TZolhNLn7QwHh/HrGgBK0/gao9Hl
34ywmXLWRgloLAAA9SvRj5VIBZQ7DFE/gbF/eZPYyWBJIWamOAFd9BCTn+fya8Oaf33smt16amrk
6wJy/N6hqbYSVDe27rNvN1FuoFRNyIpINuSmHGXYa+82hUlsNwxtpqzQK20g7hu6q3b6LmZrR9/t
UcDr/gMHrFav1bvyl4QxS34KxgtgiL1bpy7soZOAqlwI/dXhuKxljR0S4DGpVjxfn1RoVblSMi07
hs86qK5re5i0zbZFI59T22A+XmqCkU6ufhWssX1b/g18ParoTwyivlq1LI/hn6MlcjlArAl+Y2y8
SOJjzKIVy8CD+obqIU+znk9VpqDYBEdelq3s6Zbs06gXiWLng0SnedtoYLBV1OHGn+gYbATafWFe
SIgrZoG8lJ0+10BxEHHH9HmjCHIvEOTznepppcdyQZjv4iNUjynQiZSyUwEBOK1jPMvsJOAf/RR+
wYxuM183BBHqBPSEVGw+9ajmYclLbMk2TNYzIY07HQzMaqwoGW9U99w2f7BGooUJcMiMlZJdyCEm
T2IhvxJGp9P6X8LQiOuBz2U57gS87Z6DDNtweVR1D6YYhHXA59V3KG1IQ/czK6QO/A352A/SYy9k
vY+qNQqPgm0lYQoHKde/XF5E2Zmf/vrtfHTpbCwOI2IAf9040V87KUpSkKBpGJxvo3MwIL9XmKKO
Y6eXNw+1a4kgiz7PR1BtvDe7tXi9E58a9/v7BV7gCzz1Sywh1PdjlAeR7tMWOzZf43EPOXZJL9mh
mtxbUjpC8NdoL8ZLx3sZ2lWXMRZIftMW0wKUqwkVcQaqUufGszJD0IJHftjkuMd7cXbkzMFuNkbV
TU3596TWirlbjJrskTMrb/rHC8cD3EGpNxP1zvTDeP/Miv89JEwJlTaRdjkFNVZgVeZJlBuLLcpK
MYkCs0R0YQWZX19pfz/dv+Ihpb6srA/zKVRidLto6K5HtjryLygmBzqQXasjLpoXGdiycbqb8udN
8zeTwJx8IhC1Op1Rk+Wg6CH21bB5PdatQ6SLy2Wlvt7egIN/8FvIHA+Kgp7c8wRrytHkJ2OPbQp6
/Sxme40Avsb+Ea/ezRU/3/RBkge8VgLA7/13yYp9Sdg2SYaKcAZ0KxwvEuKGdKLKPZUFOM3yklYT
R0++Eoh3g4g1PVMHVPaSY5JSB0lZmjN+cMzRi9lBmKFUJS50ewjB9xncGI3O+0DdFFMClQD32xwM
5dt21KWiGcc7wPdap1F5I3ecg5QpXLtMz6IHQ9pCLH4kcsKNRGnS2t6FwQsXez3dsX4fRK2ln39S
GrY9ndVbk8yYUwd0G6ghGSAUfviYa8bBkDqqnlIcSWxtM49vfdV90VQWndHsE5kboUy23KMWPWG6
OwXu9fTVwBGPuKeLOh4bgTE/63iX9YBjcU0i4/igP6bJUavHt/wmzIzEUBc5DAFGUBV/ocgq9xQE
8vnUmAnenxz0/TovIoPIgYFSt1SrjA97ISqyG2ghHYndDImAOU1YLFCYShZ1qBjrqhO/RjcVOBgT
Y5mipgbReeSmje8ZXRNN63Z7dWfLFyPhiOuZSVE1NO+0+vvFtcNdTFoeC76PnJgXecVPLTyBC3ja
PDHhtHehjb6OXvygjo7QHHLYdsZrgzydCjEorEQLeuN4rKTTVKvz+eB1NGOx1SeGBerAJkWOPhS8
+H/r6KSekm7q9yBzL4BRWMuG64CklbOD29yubmS1lzKUxguHd1excBXhrXzVSqYW3LMwKfb8DqMH
ib9q7wnQ0a9i5yxVQA805PhIgxW3cV69PtFO5k8Cgt6mIdJH6j85tm9UoKUvoJN+3c0j/71NZDAj
cuH8rAoC3o50RXvILH1AqJwpg/6Xt0pGTZz5nhlpVOwNghi/hfNzoPeTEq3HY0J9BMV3ooKFeFNc
9hJtqPePRoQnsRgU+jSAVDkPEr232fOdcArwpWf8X1NXQUE5IB22m3fpFPspng0uBhPtevx9hj2C
8vcXx7WLwrVL8RxW29ud+9eVZPbT/Qd6DJGeuKvynv9lT+8wDdUJOGloA76k6Pn8jPAerRpxofVN
Fos0OE6xKlg8rvdBQtLBHcoaGJnVqichrU55K2r4xWiqRdJ3RvofSIOFiiuM01/Bfc/2WARRGEz+
wvOCbosl5W117yAzEHhjOWJ99ZGpyApXkjo5Gcw/erbHfSHQzqprZAzjWVwL2VGas800F5nOVeR7
Q1n3we07vbZt/Mjx+Hg49Gtft1k2r8eMM5XkXoeWNteVpWLUn343swGq3OXw9KQVIgt/BJuBtXx5
cVxZlN91vca+b5gNKMFtPniOLKUSBPLqoT8qcMbxQOI22dUw/d2IqyCfb+sc2k9EfqNSEz20HL3J
1Fo7dtmw8Y5Mx5QBXz8fbBKERIwE/IGHSEL1AZV/2QfYlz+BOkO36oDv+lZmLIsqUlD85aCjz3UD
9Y8of6jzvlcHQmfrH5zjMJGa3Rrb8UNdngzEKEXyBpMUHSAXn/KxzdzicOm1ELvXIXXbqrzX/tjs
c6ajUK9poxPTN3QgI1JNm2ANAXoIjHDEoeYxQ8HKqN/6BB6uiha3movuCvuU29spPwjeX+beKrwH
4CVBMNyOMug8zRzLHHzI0GsEw/6hFlGXhOoyaJL6kdFSUplHc+rdfQwvqMv+UfGLA4MpUMgxTu+I
NukHqnXjelFSBKpN6N6aPqIKOAb5THyw5GOt0NTeWa04Isrw8eWJ+YkcRncb+gsA06j3DpsT1Rs9
8NJ2NfwtP3wbLK2M0JIc4jCOV7DgWof2WW/UWRXjHVZ35jB8RSUzL7oRTDq/HVmvE6xJn5SEEhww
fhwQRYzrkqpDJdHgsEgvOVeSrzZgU4oxabMgCXf+LCVvQuHAX8urShleNXOZd7l+rsbTZzHNKAjH
sf2NoIaEG7I3SMUVvSLTirBZozAGZW+Z8yOHL2yU2Fd/6sgbDk42+FiT6D3hE76KJcl4IUSXKYfJ
EH+AN8pgCrKpjThijkipzMJFsRbf4zC00DigeqISJZsdCoqqmcOzRzmIYwUjXDAVCGRZyNUbSX/Z
3wlohNY4KJC+1VuxnP9e9kjMoaBFa8eyUHtyy+bTG+bjO6zBBiNMjxAUL+VSRwPyVMlY1xbecoM2
mrenJYmMaqwTz8CoP2BFzYFWttzOvJJ1qyG7Qao4gRMiXn0AkoCHNQSF59t5klHyEKZRCgSktF5k
wE0mn1bDksPhKXpzyOwvqAFRc4eOiQpnR/TkB+9UrlEP1YHtSBQY80qhxf1wkUfGtp6hKAstXKw5
jmY80hJBTN0UOdFzXa7ZJe+MEzeP9BL3A7qlkicagSCZQIKWiM6aLIFgMhKL2oPNCXJC7MRGh6Ee
Iun6dlwyqGISURIa6rpC/ZCukZyA+t+5WiKU39v598Z2B1S9sX4zv9zKoPgRBGnqDHHlA5JlGzhO
338pBhoK9qFTtTM2511DzaCLtKENK6XgytL9VdbQU0KLpaEvA5SlWrn+OQQ3dRA8NwXuHCaX+4T/
cA9xpfjKjyfpsn5mSI5CNJtU6q5fX8DnsOW8XO/D0IKTz2+msuLBuWoA5mqEo5Sobu7vwR3qjfSx
Wv5HUbbH8yHkP4P1EhyRaSsFDNVnXxq+DqPWuUk2/yco97wfAw5N3YJa1wxtwzBJzNH7KFcAYBLr
g8wGFAvg97mVpan7FfmpAIAojZ0b/0kH5hJZdO5DH+kj121HWTT3jatpGprU1WDfXXSYT0n2TcL1
8WPYKMMkuG0qfdptwCm8XoNIh+QoQMvKjJJkP2h96T+Z9sfOyBm2S+xsbQK/ROodyoSi6hCG6eLW
r56+PIXc8qOOwr1vvNZ67sdRQryOlyg1faKSlpQSP0BJXbjogwuUSKUoGPo4BA3EmclxjpQA/5fH
PghH+wJOrF2wAerPGWRt/CJnNt1wCSCteGKZPxaZEBNVKMQvHhHOCqAz5QMCSjUz7EPD8DmGT+MI
LBmzQQpWXeSO0O+hKZUeR4t9a2zyMOqTB8FgWMafkEo7PyElLqcwjy1UJfSGUMgvL4osB2vKDoSu
wbsat0iR96Rwre3UaoSaGMsMMCZWK+AoZLrr1e171qza63LWUKZz9mrSF9GYuGDbOEgCahOByeMO
mMG7hc367ILQo2Yv6HEtrt4+CxpuRj+qWJbf9JQFt+6qvNU2eBzgHsKG5oryw/ZAn5SMgL/fPJOP
5zslxecuZbzuVc6uroemn5RuX4dIHKLQdP4eKgXwyzYZxRjbV9wy3+4jyMoVfj/kR3cc1IT7YnZJ
ZJTAxS9rid4JMyaYHZH9xqEL7qGsdgpwgWmHScFnJ1JKscfPrrxG9wm52xseT5keZ6zCkhR1ezBx
f35pxj5L0VuVMyaCv79bEVB93T/WzLtHflf9/Urg4DRISKqTBfnP0M4PUKXVttnuT4K/TVDXCW/E
8wVp9Ukc+zhp3KH3LqPx3kY3I4E1ZA3A1oNFYQsvcoutrgMGOYVQruOX6c6I8/w3F4ZaV//QFMNw
tcpQa/bflCWuzIArugYytEdK6USii3g75dNAXHadj0r3tAqpxMOeK1ZA6Bj37NNw3Xk8OcL/atF8
t+q8dk65ZORGuque6zyH6vOV9SNKb/3y9OOxqykaPHLUCRG8uBiDOHX5VVKv/cW41bi2vWFBtw8O
kpUflBOyXIePexAdbQNQKpnx0gHaI8LYufBEKp/490mVDyH8t2hiRYNfGks5osPkY3WOcwgTIsYQ
0Nwh5h8AHsGv11oNey4nAGbA4xYJxj0CMsBFY0agYZXdc1Sa9erA1QnrakNa8Ozqx6o+OPW7Z0lm
2d6lDfCbVODqx4M24DjnXaKPSurmNL1SCJQZEkPl2psCnMS9ftiRF5MirM5/gRPRXLUfiP6BBpZ8
j4beCOS90YLbWMT7DpQpXqWFYl1rWEfns2U8rC4x9yW8a8fDcGbaK5lnYCAdUKSU/ItgIh1eSRim
WuzrRC6zspd1nzjiPm2PTYeGsXqq6wUyR1DRf5HYfArVLXHtu+tA44CD8px4/ieNogC+qP9UbP7X
xub5NtB5nsL5Mdi7uOXAW2HnipbsA0omDKlwWftp2KqQnqKJw1zZYU8qv6ea0XTK453ELqFTpMtq
8vNdc2z1gONsQt9lqxTb0D+SanQTz4u4B3wEERmT9yNfJNC8toeP3AZx4+FUoIN+mU+N/pDHCbEq
RHvijQCWryPahDsCMeoKxoUEAKuYgMQMze0RTr6RXyQlMftC6WcqTaioXhacVjSbGnAP1NbFv2pq
9mf0QJ0gUoOAe91qIRKvrMecgu1jR2cmh2IN6dGJ7Re6HdVGIjoMQkzmn2gKr7l6YmVGMhJcA5hO
aDtkgmKaPxahw8K/GUyduw38wF6UhqfywDMB3nqy8eMOINjFwMZqSz6NaZgiVuskqCAiJrSuk4dn
0NE2bJOGx9/meg7lHMqh/Bg8l8Yd8t6vh6dxZ+R3zoXqudOWw7e2dGu6tfikuyGW5qIbwDrkDuKO
6hMxofuduHI4FQ3oilbC6CMGaMKFc4zcMUPBOyYp03LS+zPHAbqkDiR3M/nYh9HPK63o96lYGNDd
seNmA8x3+OkQfSrLCfeOGAMqY9AmtzXZ7P47NQHF2xzC4VnzEd+a2/8jWQr63cyxJ6/Xa083WPIt
LJft1NR2oP7Nxxe9ri2lEBABfZMYW8HTlQd/pRqG7ZCeAOpMs/J9HSYKil7Pz8PYI3yNHXqoHB5Y
k4PcCowG1mbqC2GdMhxf3JiY4eUPsquo97DySpDuCHg8gNB15m1h5TcxewLF47399A+8nSMpyxx4
8AUatN+I4fSP54ucLfkYr5mNiKZCBKMOtj6tlJMSciqzS8ndRgvph35+v7rdzYc/VGAJbNXeemNq
XuR2NsWd0OSomIuSq/0mCDt+NN9R7vnrakOoWlRy9ma4DbbZ1YZ9FYKjVOg/jJOI13mgmGragVtk
oeUO9boh6eQBYsjGSKmIAD5jI09nOkNODFjRVh3JAX5vQZ8tsQlCqxO0Fc9yZ+WDLg8su2QSN+v5
9Qjjg4jlQmsFU5OcZrK24//siWVGEzrb+rbeG2TK8yUnE4BaDTu9WHw++OWfT1p19CWH5WaEcTVO
tjxrjB7Wk+fwrkzZTmdy3I9zI13SzeC6+/N2tXHqRJY/LS+/Lrs7g1ksZipLVDmQ+HZAtaWK46Qw
XMDSXy/B6oHFRDvQ/snJaQleckQyQTTeJD3r9uORN8PYufbUarnBauRaHF0oa8EPrTcNb5uNJU53
VHZC/bJHPVYqz375WjLbO2LzGQM6RCGnm/UV6GfNtx8b3y9dlt7Idpn3z5yubz0NnIcr3fXXw+q3
/em/98Gof2ne9LUXiox00EBFm4f2op8fTBqynSytb79TmSTlJAymSL6SQ2ZsXemVzbDfaQneVl1g
sNDwjfKf2uXBgembUiXi0VBm1YTB2D7aYmaJJ3EP1Qdfh8BjRydyQhCtSa3hV0ZjG8c89gFmmQ9t
F6A//vSHjlUbr3jifVoDWKshcVxn3VPyQQ1a0jcFT/sKmD2XRI251JPEbxC2JTwSj4Fql2tN1ddf
qGdwl0SLbrO9LaSUl58g+8LSME/63eJdEJMqcRZ1itGkh3t4BBRjutPFQqBKRlQNu7/xSZr7Qbv8
bv4Pj83Ct7D7kfsiYuPrUoQbtCScvk2zNtxs97x9KU9D/vPBNo/IVN8nIWCMAzdoQLHpQzNJF/fM
TxpdPjoC2zCO4O1MM+GTXB7UMiRioDaaWZ7/wsFDgIewvf1JiMyWAm9QLpk6k4Ct9fvtvp5+5hja
wPcmYUNpn3fMd9Qy8QN7FDYO28N0qNSECV9XjqNfKWvvkty7/ATYNr0G0OcLBZVT+kRESrjvfs2+
XKCqevyZ5d+loqkLqQvesMPS/k09kiw0nYlIzVG44JA+eeXR04q2N1CwR5wa5HxkDAY1cH4mRQKy
rnM2jIZX408f5GE+HIoYJod/QmTjzwsZfDVUZ7r7VYFHzYirJqgYUlAv0Sn1ObylDl0GrEslhqlJ
rH6Cxxik06fp8Wiv0CzQRSyIo7G+JqjA3y7wmwi9bxReGzdIO+wxkGzAg1A4ozXx9j7MglNanXBJ
CT8ojsDOGPjKQ7rORq0g9h2TwSmDBf2I7HAV909v+YvSbyfD+CyPs3ylgBWIjymBSrDeATjknufA
yrzLx7vW7BUg5qy+HxhbJ0cer0i8/5P9lZDRl9NlbjQlR8YAUFn8HiOu0544J3zKzRAZQzJjq/8O
fSCKJwQwcxDNJUsoPfZGUt9TExzARJDXYt8AEbvXwKPwxzWW5HnwYH91EyNKqCM+b+g/z/P0Yur/
p6xeFYtl5xOQxK2hkC76+RMjtmKJwdsSXa/J8ilY8+V/N5djwTVA70Jb0LDkQxuM6Dem1j2Ypip2
ka2jKs8jSWCcIyfcvx4PK7W1GgJDlIRdO4LZncayUTz7ypl8Ja2wPFjbujIIMpq4OhqFQHP3bpR/
Olj151Xo6Oei4VH/yb/Ub81PfLeTd3I1AG1anGv8JrEPkOQ04Tof7S+2UFYh19O/NpSuHjbjtlO2
AEe33crVLPQifm/+0amcKfDL+RD4ob6aO2TlTrmW+saxgn0PY1kROtcIPxBEwIIQUwi58pig9Gg+
rDJYkiBLZgcFAOeLS/5Zdt9RcPc5AUzBCAgzSuYf+QmgkhfYTuzKNsqZlD7GgY7SmkV6Nw1BkUfA
Q8Vx3VksRv8rb+yFkkfN1aNDwTbQQLRh//saM/kDgdgrr9DRNTYef+0yvoOm8vlfOA3rcScv3G47
quU/Z7zjN0FLfLIcfy8W0VtIYtNhd1DsCxEMmW7QLvZ7VR8eBepdrz0gl/nxnaTSUjL13z6IE+SR
Jr4A/IOYtoRXAFp20Nv58nD/aqNMxyDBH6Dq3tFctMgDlb7fNsPdWuD19iLAcX94SC5C37+dr5t2
9xVTq5Wfpiky2j5RCVK9TDFYtXjPGg//KBK7c6AyEBV6rGv9HfRC/Va/lqHQroHqWk0bBtXoMlR6
k1LsSHcXLSOAvCV9BzfGVlh5f6wyc+Iff0AgCJAgaO1RseonnP6No+c4i5AWPgwmCkPkiGTsowCu
QRpcGlTFb2ZPkFUxU+cNB1jLTTw016Fr1aRZZ0caVa5X/m9pajA/WXXrtvnnBjwVXO9atNB5jtLu
Sn2Y1FymVdPuX9DNaII/C/F8m8+xpRw6WFVOp0OsJSrg13JBPLaowU1XMCPLn9vtBnWE0gJobjv7
/SmIJPmatPmHxIlau04eeJI+d6tlzj4Z/AGktUZxef5rhYhSWqoeqRGHBvxlwwGtTVWC26zrHZzZ
/tuUYgfGSJbN8UV01VjcN45gTvR8xupe4V0In9SKTfvXPlUjXGda44MKLX2XqK7uaOtiL6HFrAdw
SoAll3ZUo8GvPhTTKB4Wu55O/nB49EJLuOF52gu4NHXX6PNNWyNFGrVPvsMvmRxWSkj/dfK5gaWw
kR14qy/EoVfSAnZpGIEeRa0gGQ4FUT3ezmyrOy+/ljxBqRmTpe/OSB5z2iB/xsTlUBclnnGY7H5H
LB4yVG7MK0oGbE6/y8K7kk6D1LC9xQAEECPf2U6/S25+nP+Zhv4zbxD8XCTIcuwASSsW/JgBTQ1c
dNomSGnslE91RPlCVXsqqORbly33M/B4Rot8OqBr+0+aWGByVAowgO0u/jGinr4Ul1iO5Ax4EFgD
UgzVA9xBOJRkcUMgkVZicpkHdJOmSnbH6c3IBhTrQurRQsMU48IEacIKSD1q0t6DPMPL+24exybd
xVqlLu/4YkM4c4zHGVqBvkD1s/EMyREDWQ2YbOcVHA5gbvR2dSHdVVLjzoW0WxdxwDhEgdSkgGiw
T8x8fsKcweFxEFUVJLOC1gkUvkYUwHPIFl1QVf9E/AwEmTX7cEVsqFPp1BpCIHjTGFviWILw3Egz
fhwFOoCfgtnJlLGzN7nLCxkwMxGeGcammxE0AB5HI3QKPznh85KBi8NSP2GQ0WdmKmzRUKKI3BTj
nfnpozIQAdT/n6EG+5KWRwe9FY7yID6KZo9MKRF+dHNqGkfgAYCFK7p6GvorSLd3/3fE2/28KYDz
lb+BShNQVcpqem2kEWT3Z3T310qd3rGCswwJy/ucC9phvFKAXLVJuUU2+voQnxpCrHRNmP1hj2E/
I9ddtdbMNx2i/8MI/QIOWOZYamewq2sgl0E15+XNuTV9CCItd8IJePsP8dnQxwixMAZ5zjR4Gc0Q
sBGmzkjCN6StwI0gnNFXbxp4kzOv+1ne2dW2n+x0eY4ucIYeJq6MPOyvK0WxKGndaJUVVv0+YY+C
bky336u2hHTSF4dYJAf2aVdyNW9IWVJy5A45h9wicEN9LKlHISSoJqmlw/5GHh1d+FqL14ZRT8A7
qwdbvEmxmt/U+kM5Snpy+lHzeIoP5a5i31FWq2/bVIHBQUuYFF9ZpY08ESkY00mtPPHLsr5VvLrR
koRVyckv9g9LX1lbGHS0tZxQ9Dxvy7Em+qdByRDuJibbiaHvkZVTT/yo5mfndI/+tzJx2IM8uCtU
ynsVFChCK3AeuDQDFowj5pK4FPd4Mkjz7hXohS8AQ8ItzWgN6q4iv/hCXnq497dF/IxTTjaw3M53
CZMdgG/zycHgg5cpIUcIp3OqMc3erMrZBmzson9M0AYvgCUnIJiBp7uHXvU9Z7uSjHF3luqkSjhp
RayZE0t6fIkpATXYdzMgjch1mtaWWidir9ms3BxyGmOORZ/StAQPGkXbuW3LbzcC88XmJhtEddJv
KfVXYgg4pnGpFxBfHJYUbs9MMjsVbRfj+QUYPn8Otzh0+HWAFdZ0o9IYPFXkXdx2Td4pCzO+AUuB
zbKQlqYZXiKdVM5ngtUmQ/E0HZE7WlP/tR3v5DPe2phLsmhJ6wKkkZ0IVH/sU2tzGN2ultpnyEpc
CV/sMRIk01O6dNpZAZtvaLnRQV9WesB2DbSqmchMj4Gtuplkk7VZyX3oGGBwyA3n6UMe9q+X/okF
QeofpKUSgqCwtwHZRv4rkxQijLVeCdKKdjvk/d5u6Avp4m/W9yTHrqL6tYExlX7GjtS41NIR3Apj
LYC16+HYjZzXDrpCj4qBG1GVbjf24UMMVAvyZQ9sbdc7TGBdMFpmxvfn1VAQ1ro5z3fTGkeIva2D
TqA+mWz7jI8GsPPy+CY25T/g+rTO3/YNqnrVY/RUCyt4qxj5GpkbGnBfd27QcNSk0O1g6unLz6Bo
mOyJ6XKWUGUQ0yDcMUEnsTjci+Jvpqh4hZ2JdYHozSkIwLtqMD067uoKPsHDCm59bTzzwlLYJ5n3
55gn9BP7yxygTVSx8bPC/lB7S8wDvdeH6UFNsbjoO9n1zptBas7MPVfOTvjT6XjkeVaRV87mgk34
58nVg6yNYaf4m3p6emSdavBtf/1NePOvIy3K7ZbHGlSQIno9Wu2pHqBMWcp+LGlXWso8teJu12uG
WtmkbzRRrWU36cKd2oEBLEOWPIZQnIH9UPkhkPU01h4e8h96TcBqS6ac8Juv//jsfwVqwZaFWebc
44xi456tFcM3EHfuvw3qfBxMPubucjk7BqL9rlQvXQLd4Lirapkw+ThvbtBDyipR2kqvNVGQrXia
u1ES6EQ3/nHyTzDj5C/DS4ZZ600tl78pdyUGA76nt2md8bPAqPHcTnTpyIyHeJzAj471mZadtxlW
OWmnXsitl+PX2QZpO7ZrdNZ8otTOiTRUV6aLtigcAlczQuWtQ2UFJh8sr3AVgGY2YGHbDbpkk7hZ
1FJpkHCONm0MvKZ5kpcFcsKhG517ajOjcKdsK3pGec19kNQOQzJdyUSA+U2mti1zd9nH+vNPRFZ0
rdJyfSvefsfC8MTlZ0/tsIY+0a7LtLF5IIyRLE6/z7JmrBTNYd0L/daYkreSqzLj5JMdeYIrHmt4
CeXke4Lksn+TwoePslRxt8BV79Y9On8q1JaQ0/IIvyHQH5jvBe6bIkIcDdgzVjS14Dqqllfqv7tU
osd1u34NZefvnsMAo1IoWqdC/o6Js+xkd0QvlgLv6M8rVKtq5dnAHsXt6rZOvWHlndOnwioPqNyx
UMfDfB0xTRBgnEb9sIoo0v9YVl95ovR3++fvwycRpYVSRtciO3hJlVvhAoAsffYsV51eKFjId3ao
PB5FA87ibE/oraOEfi0Z3c0nd0euMnXZJ7gyZBo1qiqaf9uRPhQyP/dfN1L3nkTTkUtUcX+IC8KO
HmNlLXfeovRFLjomyjf5fDk8pndOPW3QUxn4tCY/XFH9ly19eC3/aYFZEQpj8bOcqAz3tbAAcG8I
KEXekSbY8veQ4SLwkk5GyO+M3BXcNXbxHvHMyMXsgbxxK44Ypu96Nz2K86khArTE3NTwlA3wjLUl
Xsy0kmdgIosvqNWprU2KUC9Zc5lhojF5FuuQTTrxZQLKzIOC/8q5MBtyqeSryOWAxC4JPogLl9V3
NnPfaLAPMoCX6uLAloZ8q5SSUjEtliOYxryGp7aDdYK8+A9J9jl+74cAvfL0vPl4YhQ9g8X3uRf8
pcvnHMzjBebUKFlolzkC5/CJMCL83OKlgYnSsHgZLapg+YT9FzT6cGyTLjKQGVOppUAE8vdWBpsd
ITx3Y/axLNNgE1LXEIwXSp8VjcazyMr+3s9mHEwjWPudD2c6/knafpi2yyS8zTGW6iI1c2W4SU3x
0tsWlee1rwOQ7JTyBa0tu8bBr9B1OudnvAHv/6jU03ZlVxSnaXDHi7Qw6Y342qJp6SCHG+C0EYsw
m1Ab2fRV4vgPNej5sc5Atog33fiGa6yxmG64tAoBljkUW4TFCdPf/plNcBJfXBnn3c+/95+Qqmke
i+oS5f9l0VPEKzqGfSxkjftq6BkexOhfoC4+i9pNakP5tG/2M+Th2v4aaedvxCtgj7yfGiKnXDFf
prlo8W1ABXnQae1NM3S0tkJkjBKCFvDgE+01LPMqLnbbQMkEGeGWcExJuuynycOx666hZsJwTV27
QZ7+3Jm+cs6rL8nZ5ba2bKpHQrZc6rpTDFSbJKk4RSMmCbxr9RBKoQAV/pJNsplIm0cRMkDALZc2
0PFPRhCPEioTyYDmJ3tixI+vJQIzBluKO/pbLdkCuVQGXJgPpw0jbF3+FdR4WNuMiV+p06FZaS2U
kGpiUw3wPTSmjJqvl0QEdkvLDwf6uZd9OYO7C6+C++FCDIeDdIvmpWDifrpNuXexnCADqYjg++vV
6Q8H/gUu/tpdGmD+ewU3tuGPzd7qnsV6RiVQkrnZ1PaHLSyqXX65F/a6nxy0Mrt6uerWiFl1f0I1
rN5QxteWRBVkwEIsSq8lra8Qwwd+Im93ecQ8XA3v9mHp5jZbv2osu57ZQIDDFaDR/nL/tAKhvqof
FUcvOeYj1C89zCcEnnsp7l59xRR6ZC+/MjubVPuTYz7khNTIGP1eJ25MqoWxOycnGkvKXLe2fOXL
uGccYqULwspnwzzMxhordyqteppQqS7mNkcwfYhQoLd2Iw+r5ejryDkEF01IfXvb2ihe/iukz0BX
SuWXCxz0jW+Y/Hk49iJW+VRvzWRfSk8nWv0JP8m/50ynkHrgMIgVY6xhmhqyC54ZOs6zA9Myicqx
FvSlPN/6HqNU7avygIr2lJPMfxfHNRIriujWo77AsVL67BBYumnxHZRcscLfUWYMblErrBmGP9bd
GjGF9jbVcTbioSpHD6Oid6qYftWgFR8GFBJfNvMBTyIkNuymEB3nu0PRHABOWcAwIF18imXKYR9L
zpxYSzvucy9O8rtJWX4+4tpMX8BVSkpJHaVzxc9D8zFrFLlDEN4khHznwrgSBupLlShTUzhf/3sy
JUqN2iON9i6tSHlSozOQqn/fCtTfQsCZCCLlVetmK5Bgdz7uXXYWj/nIBsucO7YZrFJ7w84CtrFB
7bqilxcytLitIa4tEXfnWH1bKeeQcEkJ5mDpXCrvkdjZYLIV0luY/GXIcJM1XAxI75egmYoWpN/J
7AyLCUCL2IKW9UK/iqRvEmfG7NaJ7AqarJBg0lwDygq2FLTXvw5XG9jnb109Ivd77OaF+6qrZOdK
M1lH63Faof+leozJ1yRvr8DYRIk1GiOpVU/1JyKf6lOND9t1cENmu2OP5NxZ+ECOQDl9AVa+zDjA
Y3AsvLLnJOGiSEmakCvMVA1faBjUF1YcOu14Hil0rX7qSfoKr+JEEkEDImSaZyizXLMQtcy+H2+Z
VJGS8gvmyTJQG1/pmNwxZ89w2+8JwtH22OyxnES0xbb5+JJ9U3vaHb8nJBrAfgx+Lm74nsVpTKfA
l+hJYPm05kXEtDioLkuZ5OBnDQ86zVhGT/Wt4Ir7qHYN0gwevhyCtbD0/R7itcC77w6+/EzQJfUc
e32+dJXGYv9RPBC8ZlbeTe17UxRJNYHoLXKV1YxypRBfL+8SC3g9S0Oidveyr50g1Z2Ldl4YpVaj
v4SSDQqf7PxpGHq6fsie3HHMDm4d/Byi6qCjmsCuCFflPRFGO/gjaFBnk9gYOI4dTYMJwusC9T58
j/0YSs0f2FKhCqegwa11cxklAkNPw0Z900a8oBVvVJc54kqi+q3W5+a8i60ujnsTdYOnMpriS5Mu
dUvs5uevEAK72TzvSguvGYdN62GsdmfUJ1hTUpHeBjaEe5mI9SKhPOLAVRfAriqMuBfeI0aRDCoX
3B+1YvquqShLBhW7s+pUy7CC6OZwa39Fr/+BLPGr5fmAemzLr5IN2/sDXny1so2Ok3Oo0uTlJBQm
/KEK2iv9SMPtteAAtpKKfIF/YbhC+nY8tNsGzqNmvSG/vXRPErRruHaP5inslQN7yrXKgQJ3yNik
xKGD/hHyYpWmlx/a75+lh74Ez9JF/PdGtMATZoNzsrAOegiyno4aXdbBx0m1CKi3lT2Kq+Z3vS11
14jQ8FHArt55vO8LGlWbwPcb45VDRF5qAUIvN74vv0/nNW9r6btJ1NOozsmMq1knw91Dk2/dqIhg
lGvKh2ODw/V5y7RbpXXSunSRegkjt4OmMkHTh+o9XrqdWvAHbUlqrJfLKzLQHWhVH53qZpHcWLH0
8HhFb/EjI0DRLWZUQcazsMfoHVcN+e7S9378GE1c0DtkXd0o24Jc9jzTmDyf2x+K0JB7CFSOpNON
JEce6x7Xr7YtRuRSJyMoub535TZRxZhm34099J14AkhjIPwb0c0d8CJJ5BuGStiT366VuWJku86g
YNG/u5+cCi7DZV/GGRb6s4E8z4B7a2oWQUsDSj+og8Olz1RQ1byf7sSk72IRr80Nrqd5wKOAvaR4
OaRxS2aFgD4SayrPu/L0CylmFYhY3Jo3CnyxOJWJR/tuSHUHW4fMt39MqLYL39nPi+a57lHSj3Lg
agSatf1f61lVs6Y57dA+LF/muv2KRwrMHcp2UGkquDIEiiaeMLOqY7KaQwIs5BnvQYtayF5NJm2f
l81ozcvBxcZOLRMzzzx792zd4jUoMIwVWkre1Fyi5jKoHUJAt0c6/loMxL4EV0x10OmuFfIiy0UB
4husKfTRyGyXaf2Lw/uYBoR4VLhL6D55aliewQyAL5GwhcqqAhF3MJzyyHzAaLkWzC+Ap31XbxTx
fEKpl/kUWCGE900YOFpA4ubssMUYb4MktOlmzShtnarqYFh5ABlYpnCXqTI/WmcZEspQVhKQZfWP
BqhVUFvhGZOjHFjxQ1FVB4r76gqBdNJYjp4nAh3mvK0aPNegLwxSFH7FKUe6e+LxlW8zQm3Gorg1
rI5WxckCl9+qSwDUdbtfm+iadah7MxpA/V+OXwXIWc1Y0Q2QCQFF/swDelwg/Krvhp0nu0aKpghi
N8dpyoDNuC2cjiNFPf0BbkrkIaxuYz948NXRxrD8alNVgKBI7V38r44qPIGMz+XsaxV7dXba032a
d8sLkoBG8LlZPINbveWMyxvtPWRWsVPR/+FM4Ob+dcRmblaRXMb2tZZWTOi71Vw5UN//A+QKkX5R
DUetkthc5YsKUvocd2CPMk4XjFxnmBo591hSWnzebysQk/DaIi7guJU+dBAFkPuXnGEBf4VzlA13
qud5v+H6DV0fsZCsoPknaIy7a2Dm
`pragma protect end_protected
