��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�GN�Џ	�Uڨ��ky�3w΋���Fs��)�%�s��B��r�uCۯ��R�?h�t�.�:Z���D'���c�_�<gO*��UwX�/;�P�N��<(˔�ě�m��2��Y�X��U>ҐOy))������R5������^���;k � �� �w5���^-���w^��Z�k|�Q7;b<o��?l1]G�N�L�ȭ��i�kGN����5�%�Zk��b".4���� LZa	�,S�e�J�Q��A��c�}�!w���k���M֗�;��S�[qԧ��WR�L�a� lQ� _��tqA2�l�E�Ӌg����'�/�0��k����h��x�fFd�6J-������+$��P~P��8��ng�B�l��`���iA��uS�����D�9�waV����2}Fe6��BM�U���,�F2!�?�{�u��Q�T�_c$���A���hֲ�r��w�;x/�w���?+���IP�i��9�Dh����a��V��$j�(G -)z�g�x�� Q�'RY����ks>f���n��du��(�
֢'ژo`�I�R]B?�������Xj��ꮚk��Exkn����̔!x�ɻ`u�A���{�����`l��ѝ��'�+��H�+��h�G����A���Ì6��3��BsLG4�Q�ZC�LW<s�Ϫ�nw����bF��sxc\E�J�H�z]��B�쉚�F��mCq�r�d�4bƱ�$��YG��.Y��UF��R�4t'�X�"����+y�>IQ9�AY7	5x���HR�^w��_/�T��?�	 Y�|�u{͟����L$r>ɜ^gE��P8X���ܖ����HTK4�R'�zh���l�TP�/��o��h��y��)�5�$=�F�~��Uesz<9�2��*��0�5G���2J��p�aƆ��'�ի��\�,�(��>7�y��e�jD�<՞|:&ft������e�C���5b,̭�&ƅK��m���`�Sm`�}H��T?�^I��AHC{�cN�_�E�
	�N��gv��Q������i(�=Ϛpއ<�w=��4z����� ;U��}(�4�CY ��#���z��J$�fa�[����.�Q>�>+6��օ�V���zUF���7�Jz �U���g�"Y�YQ�CJ����n-y�m�1�'Ϸ���:c{�ݡUı��L�D�����W�w���3�~�mX�RbU���Z�rX��ty��7�$T c?8h��hOx���if8�7�乆0�YX����s m��<�4�S
���3HoplK/�����o�k���7�?���Dt�쿚��F����-�1O�<���Z����c�����O^<[w{�z��mWp�Ap ���1��5������ ���E����o;X��U��m (���Z�p[u��"��|\�'k�/��),�?����ey�=�$"��osw��h�|y�G�ʢ���Z�嘏�?����u�!� �=#O�;�қ	�MD�Z��'@>˩� ���Y��h�v�ߞ�Ia�Q.�S��)8Ϝ �h�Co����s�$/J�
�D'/tR���WK|�u�����G�v���t�Ȩ3�
E����#;�@�'(�j�4� t$�����(1���h
{h(|��1v�M?v,�T -������S��\}���,�)��4}�� ��Ǐ�3���zs��O� �L'V]�S=5C6&����c�/�~�m����!@g��QOT5H�������c?��?���+��Ln�,/�F�Q��
��]�n�v�h<@��I�硟���pf�J�9�W�=.
�M';���{BFQo���͹\�Lc^�����x��7l����ٿ��D��@���hk��3�����1h5�!���&�s���T�Ϫ9��1���)��}A��d&3Ԑ
�����B�F}�B�g�yLzHE�m�zGq��;���`����-��y(��d@1G��{��V���\	S'E܊Ie�oA�'='��Jv��;tX�h�������*�Q�ʙw
�e��8^:����jd�\-�(���K~@�BG@,.S,��~&� U�2w��-�UzZ�a�x)�G�_�	��4#����grzi܏�ƫJ�i�ҧ��X��r��9R`k�l4�ru��㤘�7!ʨ�٧�#<�QFȓ����YG��usI�O�,�v�[\��93f�%�	 *7�0K�����c�O���3q�iqT�O]*���&zd:PJ@:V�v�(�^�5]'�m"�仠 6y�_H�H�����b5��%B�S������TW�{�N��vLl�d=�@Dz���K�^?7t��{ׯ��!�WƎ�` _9(w��LE�i���nC���j$�3&_��/�؛i��`fF+�����$A�͏|����k։�����̠b��}Wx`���_�F b&f$�����Xk��g�h�u�(ŵ�x�w�ϭQa6�?=a�Ȑު��*Nu/�(#Sl�+7�IAk���!�t61�c���36��1��-%ud��>����/��챽c�$�Yۘe�|!m	M��B�^j��N���q�;��դ!%�ܚ5<{/)j�l��̪�$��.����)��˽M�x���4'1@ǽ�%1��"��I󮾜d5�dD8q����U��]��V�!++?	�71^�g��%⠶zYR��*l oP!�F�}�,q�� �\���=���E[��c�Z�Ws�A`�ZX��X\
0G��d�Z���f��O*;?]����ӈ6���re�&X>_E����@��S%��2��K�O���g`�j9w!s�^b�Gr�?�-��e�dYg9�>����ߍ�i���?5�Dɓ��������ǽ��`7ʕ "�����Na���Mb���9^ly�1]�Y���g-ݦ���ٗ4E���U�}6��h/��SW�Tۭ2��OS�6���Å�J�CZ��x���4�^�-��h�ʕ@�V��\��������&_I�\^�1"��υ�tʚ8�_�q� �,I��if�~
�����C+tEZ<��>:�{1bDs���,0;.�5�R��$z;��h頒Y<�XJ	��'3�����W���"�=�f�!^]�@ۓ������15�ᔑ7�Z6,T���d�LS��&�4��J>�V׀��=� �V][C���������_}Ԣ �v�����%Y:�~��T�Q�+��j~�KI���<x0��%#�3,r{z����&��$j������%�F������B�VF%�qє�Ef>��j�}��<��v�4쏽>r�%"�9
�O7y�vH��=�B�>M(� �]9.W�P�;U�	�����4�(�l�%���o�場�<ǡK��p�H��S=l��
ܠVd��=�^�4P����r�Ɲt_��	��)*�}Pk��߶b�{t���WRVT����/nzS4�-0쐠�bſ��?RF�R�^�woYms���a^��!hE���1�59yI�f��	3��l��TirH����c[���Rc[3w驽�Ώ�i<��!5c� E�mБ�:��ެ���37��FG���9 ���p@���TZ{��!���`ȃH�<���"�?DK�c
$	�����y�Y�7������)@�$�M<#�4�^�����)�j�� ؉��&*���ۧH�=���n~�ۧHMİM����D�1f�����oYʸ�}}W_]Zc\��RL�XQ�h�M�Y�@�s�g�b]�9�7TJ�i�ܘ�I%'�"��(� 6��+p?GWTI�)'쾌Z���HH)�3��qd14��k��I�e��.����r��. ���V�D���K��.�
-��SuO3�m��|�ȋt���(	_�U�:���^�Ň��N�v���{��fQ��ìb�.��&�i\�e�*��.���se�pn���8n��#f"`���=\�������8Z@���|���xw=l���6��vU�EgP�͢nc���g������C�b�f�m��LhO~�����K�09������'D��?�f� WnK����oN�ʌ���A"� wq��©fc~0����iD���r{)�v3���A�U7�j������g7�al�0s;L ��"������v1�t�uQ(`�o�|l �o�cXw��/�=�Y��nt��F���ҤgL^�����"/?�mc%��S*�����@�>uz��Mpi.pENp��m����p�._�<|��w6���|W
XUpM3r+qK��S���V�3��p��p�JW���hU�,�Ւ�ԵG���a�����(� �2�@8Q����}�*�{����$�\_���N���cf[~��%�5���\7uk���߷䦑.�āM�h��&�8�w�Z ��L��[���$�����P'{�V�~#�X�@�T'ss��#f|4�vT�<$�ֲ����L�Q-�*���$�H��*��0�\>3���H�rTʙhھ����	o�!�zk���6�?����J[�AxR���*�S-fVD�����}�=֎D��I�l�,�,�����Y�ɠ���ߺE��O�[�σ�����Z����(���*g��E�U�h�O�W!�>��d�n��-c~ӯ͑�1̀�v�P��exM�k�����,Ͷ4�R�j2��o1�#�zg�� ���\϶N���͚z�w�ДPaC�z���V�yl]�ɓf�y>,wF�C�=9D����
�Q�|����3�5��'h��jVD��� ��� 	�'g���)���8%�Pvڝ�RA��ɰ���f���q\�0��d��:�/kD�[Yp�#���*��?:<m��8�L�{H��VИ�ʕ���@$r�8�SP���Ŕ^n�\};�ӯsL��^����ׯU��Vj�W��e� ��>O6M�"�?C�!����ڑ~�c��%ΛT����>�eԒS���W����2'�QL֐ˎ�quk�ky�9ݹ�|���3��r�襍���=���۟m��`Q ����Tg^�Q���ˮoxg*E��R��
rF6��[��2AK�8���| o���A��K����h�K�~/Hˆxu?�&=߇gu)ؽ���@a���[}d��u�<;�.�C}"���(~5.)�EQGÞ�M����v������#��ڢ���Ϣo�TMg9)��ȌN;f4�Q6ԉCs��3�D��aۯf��A��R6�N����6��q������C@~���/�q`����4U����j~wݘ�X.6���~�yX-����˫(2݁I.�@�ލ�k'Y��})��o�Ց�l�|�Tlo�p�`x����y��dR���6n�c���#m�k�3%�{=0G�f�Y8��a�1A"�����~�Q����a� �T!�wC~{��:���C�ۻt��0�_A`l�b%���3g�w*Q�Y��d���b!�a�C�q����,�w�x�2�+ƻ��_��S�h�P���0�8Yo�������!D�;�m�.��E�ID���Q ٴ�u�s��F��WY�����4��0v	���r�TI�a�p���}=�mD�X�Z���z��.���C��Ev�������m�9�Qr덄�u�'A��C�B�}��9�	�m
��US5ٝ�ԃ��~ׄ,���(����n����a5~��k@�c{�Sf��7PP�e�����,-��8�Fb�}n��?'��6�ZI���y��5E`Z}qit�o��!��pq��N�ft�6a,��3���p�ZG��f2i��۹�tb8��Q������M�G>�n���������\��5���H-���YQ����fS�i��
���ys^�
�4�Ϥ��-9�w���jI�k�^z����cy�l�3�~�9P�O����7-=�3@6���se���Oa���'��L�v9R��ї������t������`1�H�t��Fj��"����}���O�8aw'������&���>��!����)��6a�}�W�E�Z
5�_�~�7��k*,U�IbU�� �&�#��/���~S�����Ǩ��������\K�����G�&S���}3�=v�{�EL�_M?8��;�D(��.������q셖�^��h��ݶ3%��	U_�
1T~Lzӝ���u}E��%���"�!������J�֞|\A+)箋_�f����\L������ŵ�Ƈ�(y9]��x%dq9��¯��?$s�a�hh��8<HlWPbX��ƅ�8���]���e���ŕ��rC����Tma������B��[P�$����*��5�Ձ�	Ri�:(p�*|��׆��,���G�;��I"B
{q��E%�:��1*>�mD�)�&�sefyEj%����;q��<��4�!���`���	-�x[k]��f�8}��/��mmKU��x�|� �v�m�����X�O����ц�k���^��'Y	6\���MDg�t���nS8ι(�br��xTl��@wk�R���0�st;�Z���lVV��A|,2q�E��?	����ڱ�<��꺄 �G�^s(��)�r�!�dkep�.Y�_�0�`�^"E����,�>*(QRh=Ѹ.��	��g�U�<�'W�Uc����_��I- j����km��ԏ��
(�ȲG* ��V��%��f*�h���z�W������D�tk�z>�Q�������x �Te:�g�2��l ��xY���X�OP��م���|2w����\����&���Uȱi:�:m��ͪ���kLt����N��V=9��B�л�m�5a�����(G��?�Z���DVDDQ���i-o�����M���TU�y�塱�Kh���U<�u��-�=�3�e5-���6��*��lН;0:,���Q+��~���?�!a��1�`ao�0}t*
���0�.8��#�=�C�D�W�{��5�̊����4Y�
��L*j�5�:k����y�-
����F.��kps��[�� ֿ��I�j�rr�Yhכ�"��^o�Ю)ݥ׫��T�f���B��`�-�L�50�2���4��3b��Mqу�bĶ���j{��]��)� %.Ĉ�Ƣ�0CxvF�Q����;���e'����e	�TP�������u)��
	�ŀ�J}N8��4��s�7rl��a�'w!����YR��uf/�:]�+��}�fx�����͂�QmTt�>� ��C�Qfq��{1�)����[��#(���䠒p��.�\��q�� d�F{�MK��g�IS��ߩZ=��zyB�;����v�9��vYb���2?��:���M��n����!|9������C"�[����+3碢�Nd�i�k�8�V!���nK-i��/�l�������yJǢx��f�x�;cN�{��a�Y9�|���s�~���a"��TSF7�O�&3DҿG�c5�xQ����w��k�l�x�]GW�+�lCa!��<��B�Z�mD-�HJ���%���l�w�3���O5)���ǟW�8�,��]��]_�&�͚H%1S�S����/�n65~P%�Y�X ����ȼ���fHjċOW���i��5����)z��=;V�FKl̹�!@%��&��2�n�-ג�xY�;�}Sk]� 8�U�E<�;��7�mM»25j	�8*�J�σz�=�9 bn�����?)�8�Ϡ����%2/4#��\���VN����ѿ���Gl}��9�C(�M=��^A��®�4�_U�gyT�0��ڲ$�B��3��4��=�L/@��KЬ@p݇����c�U�M�g�[H��aN�ޚ�o
�~���:ag��zɀ��(���J�O��V���Wm�Wd����]x��q�.YL�fߩ��fZrf9H
����f7Ǎ�pEZ�/��N�	���mg�j�-�F����|��o�i�\��5�w�^�"� Sr���t���=���H�����	�R�b=8�pϟd{�f�طo�������A��h׫�G�����{��D�� ���e-Xl����h�e�}a�-�<�Yy����_�����n�P�P��(!���C�m�b`�ǌ.�+p�-螦�z@�U���8y�m��	3�OFDB��㹂�LiQ�Zʃ
|޶�%O��k:X�M�c�gT����o�����;!Ւ�˿����о�Ύ�Z���R�9��t��״̙�$���β��M@r������O@bڇ��`�c�͘eɕ�eŅ�6,��(�2g�f4U�b�������j7������s�Vo���P%m�N���G�<�7h}�6?tQ2�޹�Z��\���l_�,o�ޝ�rx%5N�Ϝ�7�C���06�U�SNDh�=�X�@)�����0��W��AM�:`?��-;%?z��u�iΧ�[���9@Z��/��2w5�/kffQ����|m3�2�]OҌ�������V␷�7���i�t=��XXXL�Ȕ�v+-h8K�R��ڈ*(�q��*ȠuB���C	�E�(���lm[.ɞ���+� ���%�r�=&�K�	{��%�I�+\�e��k�.=�R=&_���\{!S3��jo#ف��pLc���=���ܢս�ZM�������ׄEe3����} ��[eƍ�~�t�0�V,�2��	��DO�yd���@_�[e _qw�u�%J���d����<c���G�hh`u�,؟s�l�O���L9�c�U���	�qD��,�����u�1q�p�C�E����*�q��z(�:Y�ȓ6��l�SF��F�i����0V`Z�r�J�FL���gT�C2.���Į�[�9y�o����qF{������A��=��T�l�z,�C���
F��p���g$��Tю��x6��5C� ):S���K�$���M�T�TQ\0��Z��l�U�/��D�C ��)�.4]�%�~���H��IU�sF��*1��k0��������n
14γ�1,��?�"MxY�@>PXxs)��PQn�`0F�����Ll�+٠����k�Z�͏��'9���)�ݒ�[T)�@3�;�٬n0�-S�XƽY�{8�!X��BR`�����$�X��G�n��}{�{�z�����4���^8�=)���H&栶�[�ɮ�*'� ��3R��Qb	YϲU^�n����a@�����WǠ�B_񈥌[W}z'��큻Vv�>7"^�v&�G(����#$9J1{Yt~��U�j�����H�Wʊ���@wv�S��M���QiY��Q���v�SJ~n���
�j<�?�#|6{�3R'+�d�Ms�2u&H㌵@n�Z}�I:s�X��ɿ��޻� ��E٥॔��lH`�sp��W��ˈ h�A��"E��t
^���@����ֶ��V�WY��d!ŷW ��o��YxjE�.���!Nҭh���gV?.�<W�5��[w��[�/�!�.�7ž�1��ܽ�3�+�d<Pvq�tD|JJ�K�Y=�쟾��.�d?_���2�O��aP�݃�
V�ŚT~�hR�+uϋ������9�F� �L!�"��zlL��g+x��
i'�����r�����?�r~N��!V���Oh�e���D�u*u'/�||���<^�"O׾�;8�}�s!��K�R �	ǡ�0 Ӓc$M!���<B倸w��o�*B�C0�1��MR�#��w?X�0DVQM�qk�4�z{k_d/ٯԫ؞ԥr#od��>�00�X����m�-�����]_E�aTd:Ş�u:V$�O�o�ʪ��|#�&��48�=�{&�]�F����Bga�K�=/d����LV�bS7<؆��y4�����Ψ�F��iU�2[�-�П#$�T���DGؚ����d(ָ��EL'��,���^��1��ۨ�_y��S/^%*q�9 �VgC�SaȻ������yAF���W�]���ߍ��VZ"�H1 �=W�Db5PDG��""�։M���������y��K1.���<sdM��V�uU�M�K�f����9���z����iN�=�/s�ػ���Z���~�k����+��RqdA��puDBt�(�jߙ���o<3���7\U���ȈhrX�vQ�A�k�u3���s�,�]-ߥ����Ო�T����egi�x�^.����c��Ga�Z�Y��$���s&���H����k����=�A�V�=��>ۖQWo�lLH���zxI�[!�hVgi!'^��q�d�cR����_��
��&Ш&H7�Hs��a>�n��$��'��=7�#).�����4T���K�Ȳ<T�F	���1^�2���`�-�[��r�\��ZNtE�$��
0q�9f���MM�`�p�i���U��k
B��>nh'���-X��?i��kS�Ŕ:��z�l]^�&`|8�_'�d�|�����t]ƣc��������E�ˆUR�O�C$SF�E쉎/Q�AA�w`�	�2[=نzI-	
ۅ4�l����-0%��qӔ,>�?��L��4�髰J���V���VztsM3׵�+�x+�f����|�Og:�=��a߽:@E9�á�BX֎�OJ�F�&5AO���.�n܈�DC���ODk�j��֙�c&�nVP�q1�~N�T���u��w��%�iEp稱�u�Fm�P�Ah���x����"�FK!=�z�Ϸ�	Ѳ8�����C"��J��!2Wc���hbr�dc���%��w��-�P�"���4.���%��)��2 J�'��k�*eT����'���!5$cl���:�i#���@�Ay�;g�s�XL��A���Pb���U���"���
�X���F[�EL�I�?�UM��z�=���6�n���u)�j>����瘦Џ uO��m:�ŵ=���}�A� tf-)���+����2Y��L�	�\�4�ʯ������24w�]X��G�?���*.aWhL�ӿ��Uk:������7�0"CiШ�l�+VQ���Y�^�,�+n��\���x��\![Z�$N���8m��Z�;�Ԁ܊��Ohb�S�R>O}'������Bs|�I����\�@!���z���YQ�q����߾|�2x�=b�b�$�`k-n?�~nY4���(j�&1�>�ARb��Ƽ�ӫT!��i������6�o|N�������;�r��F�����:�IS���T�����,G9�B��x��5T��^K�;�3�����'jr��7����8��C	�8��FΫ�y-�Id��Ad�#�vI���*�+�Fj����^�y���[�L�a=������#7��d)��/���\3�K��4+~�|L�U�d���r�������j7�4Pˮ"5t�ן�C��Fl��B�bZ.�g�� Dz�$�_zZ�y`�P�@Ƌm���-L��ޅ�K�zjSCN����/��h�h �Y�$}�tf*�$����*�o9+�����1�� �Z�p�z���񛇤���i�mz�>�6�9T��>ܫ?O�Wm>{����1j͒y1ۓ�mb���Z�`�jgtD�jE�Ctl�KTr�\�������[L>ot�$LHXr���O0��0��#�����I�{��
>LY;����`Љ���0O����)jS	��c�+��6�#�"d���NXeN�f%R��:s��E�x)(N
}L�6|c�@�����ў%+��P7l�geN9\f��.�I�t��թ[����������+:��F�P�̗hhw�`��'��r;'�XURםl&���la}]\d1+�0ƅ�H����x���C_��tU�j
�.���ϳ��ON��f���YD���Z��9ԓ�n������m{��&�>�Ǳ#!��8i����y�Mr���47I/���_��g�N � ���X/dvT��ش�cF�{��#�oJ�'�s3YWY9�����8�]Z�ť�mb�d�m8��w�_���n����/h&����6	���:�&D8C��j!�Ϳ%8m�t��ݠW�E��i�2m"�b>OW����`�4k���3�?E����a9xf�k(�l6�7����������~'?�#yׯQ#��/�+�l�(n&t[wM�+���k�+�lʄ(�S"cI�`6�}�S3��c`3+��rx�Q�~lv(�z��oʬt��B
�Λ�M�A�7K���&�
�f�*�E��c�Z8ͻ�s��*)��1����:;o6��F��˹�(���\7O���̢�����0hE��]D�r�����ߴt��!�^s�8t P���%��|=1�SFј*ۑ:&�s��w�@�`%�mKB%���ǈ��n&/u�l�*���SE���ƞJMiB8�eN�2���I�C��P��RM��q�hf�n	���JC9�S���GYm�ýc|z2�֣� �B���V�,����#:g<&�ZA�Q�e#��V͵�6�dqd�μ>��CR3�c�����,�L�l
�2BW���w٥��h� �N������>[�Aå~�8��>��\Ê�� ��ᑣT���Ӌ��߿^��[��8}{ЂC]9	���!�d��[iX��A�6��Cq_�<
�8`�� F�����Hq\�DU�m�>���C�;�s:�?�v�yF%ex�m��ڣӧ����ţI��K1|`y��b;D���8y���>�SfM���lSm�@D3�h�>N����k[�a�l����e3�y�������`TA�3Bt9��-��� �|��ǉ}\����x��Y g���b��uy���2$���O�*:vZ�����j~-�����#u%A���C��"9���P�}��J遰����?��Tՠ?�2��5��Ư��U��R�+����&��V�FY��LO브��M�*ǅسR(���Ϝ9a �>%l��.GB$Cr�%�D&� 5����*�vJ�m�_���V�{E�j�S�B�r��ڎ�v[�����MU��6 c�ʂ쪷�}X[��H��/�i��
�~s6��ٸl�Wh]C���W�	��թU��J����J����U?Z,�d��Yh�e2Z�!����sM�˂2���Z �8x�Q<�_v@�<�#�a]��;�jg2����\a�I�Rt�2hG�Sƪ�x	.J��],�щ�B)c��_vg���h��9��!ucm�?��F�#n���#*�R�2X8o�N��`��,;�鷸zo?�{�t$�!�>�-�8�C%�mR��v�m���C��j "i(�ׄ��o�H�{�:���o�v�@���Ϳ.d�X��Т>K���]����'b�+�v˝�晈*�NF��6���}�ʧ�pg���i���U�*դ�~�
��V6�V������z8��u�;����#я8p9��ŹF^�'6x� �~����c�cg�7/@�����j籺�(���[ZSn�۾7m�J�/$�q�'~�+M��č`a��ႜ��
�M�J).��%�-=�8FT�|	R����}�i�*�qa�V s�(K�X�ަ�)澡�����]b�o�CjHA�3�4�Y��G�(�'	�ᴛ6��m���x'x�����YqYފE@)E�h?�U�X�S��%��6Y��ej�\��>����o* Ǿ�N!����~1JB+��Jڳ����77��$ȩ:$�iP�iF�h4�T���9�Q���� �.a��㗘����F�y�����HR��uy��V~	?�2�v�H�j�?4�р�2؊�{�j� �&A��R8	⒲D����ƴP=��(r�׀��� H[x�=Z}Y��vRN��0�W�<���Jw��ϳ>���R�я�/�
�~ o�4���j�R�e�8p���1�. �����T��9A�sH��8̼4䷑�$wɤ�����`������Yկ�0�7��t`W^ ��p��m�s�_m��D�A4g>6�B~�K�[�ɯ?���.�經OBɻ3��A�89��o�f�Q́�s�"Y��ޱ[C]Ɯw�2���&��b��"+����6���ɰ(�8\��b�q���(���5¢�����*��xcuZPʆ���\[������U���
g������*&:0�N��ZC�^�j��3>�!fՕC<���7EIl%|��:[�X$����̈́�gF�|�2p���vgu����Q'�q@��������Eg��'�
�6��OkMō%n���n����г���LK�fyq��xq�+|1<��z,�T)8F�/�&�(PJ�w�G)���ӏJB�b�D�.G �`+��w��vtzE��+�[�|�{��wUZ+:}����� J���L/N�z�x+�j���:���Fd.(B�3�_n��s��*_N`׋͓:�c����3~���!j;Nޚ�<�N��0x���ҏ�5^�,�(����j�#b�{K.Ϝۆ�.����}!u~`j��0�*����̞�pEŶ����x��}�1B�Q��E��`
,��)�v��Su��=��@�����}H���Il�O�� h��PHq}��|��z&��(��V }�y��Z˓�.Z�_�����P��Q\�'����ۚkV�g�-����<�}�����'���P�F�A�]�g�m>��X��l�@�Wf��}M!��|NIy�A������;ҩ��*�RҾ�B8m��!%��ucwՍ)�\��I���~�	wl�|E�*U*��l\�4����?�q�[�	��m���)�ѳC�ʦ�qi��h�ߊN��u�3�@�ٲ��2�,. �[�|(gh)���~��k��� ;yM�x�g�D�D<��OG���V��X��CZ��	=s>�hC���$o.���%��bt��0�p&�$�����u��쏏:QO�@��U���;$-g��+��DJ*>{4!J�3���=h���P�/c1�F|}�6I.�2F��%�2@[Ý��K�p����=�IQ�{����g�n_��%z��Π+J+9K���0�\-2z�P%�'�S�P��c���"����u�1��G����$��^BK[12P��A6� �
�7_��:sr�����`���'N��0�}�#���wĪ(e:m-m{R�HN��I֢gA�ƿO��qءi�U�byc�ms�B$��S����q�R��@�#D<5����>�l_Em<�R��[C��-�-p5q��^�R(�/��T3�i���{adqiaꟶ�fGc�̽U�#�([~�p��C6��ے/�}��ˏ�(r�,��Ql���1ܔ�O6#\t!��A��غc�T3T��<���/���<�������#�+�d��毨y�1W ����0���^Ʈ-�� �U��eȿ]
h�+�O�"q§V"H��wt,+[�e�)�V�Do�z������o(H6Kѓ���D)��М;jG�c`l#�������y�5��ޖ1��,���\�|9�8�b<�i��1��kg�_H�>��3�,��ϙP���z�����"�LP@�����S-�C$�ICD�M�^��d#���	J�5�� =�#
���`���/��gZ�O8�Ѧ7pPv���=����Rh"��¶	��W?����]
S%^g�Z�*�l�gb�E�l��{I��h�AX!�$�b�H�M�2HM���@�q�,�����Le�o��/mj��i0�	�i�-M͂D��0l�;RE�����S*��4�aF��' K�TݯUQ���}�(�s�$q#�P���e󙸹@	��l���9��a��b@e�h)x��2�|�e�'���,w�+��C~ J[��.������GU�IY�;m]֐Z��5���>
��+��R�g(�.�����Q�8Bc")���2=��fh�.������<�ye�0���=af�50�wY�6�Ā�6�2Ř�[��� .ó��[��>�qc�B��GKJ �x�����W-�/b�J����.~��Վ��'�W����r�.]�ܳ<����hH�}u$I�YS�+�;���[�0m�|�����cf���-G�|��5s�8�񗵭�#^%�بɢ�hݤ2����������$l��|�!�6r�������`���ط.���w��5Jq��C\LH�s^s}���	�;�-R������(K�� Io����+�kL�"/	s(\[mm!�����m���B�N���Z*�=T���	���u���1�!�(���!��@�C�j�t\�A�9����B�(���}"��Ʉ��
�'ۣ�Q�l＂p����PrչV C�<�a�ͮ5�Q#�(�Mrxg,VA�-�
����&ʄ�Yw�>;��\މC �Ma���ٮo$|�pLW�ܧ�����J\�{Fҡ.(��A_M�����T}B�,��h�*}XR�i�üb0��v/]�C����|j���ѥ
��ŕ9�/��m�=P����D�?,��Y���ȱ(9�˖
%���?�jd��Ui:lM h�i���ͩ�ܯm����3�܉��^�wygp⽨;.}K��1��:��԰��F�g��z?$	�v<�z�����4)y��2��|3�a������n@�_]��,��~ �Ge�5qpD�*E�w���|� �o+��$_�I\�p+��ؤ(ڼ�u�&��f7�^YL���U��@��������}��Z���a	��4+��B�+��6{�����Ťԛ�&ihq@S�}���?��!�pF�M*h�P�bMk�L�h��:�b�;Մ\��_��*�Oh�H��#��ʫP�EW��%�{8�-��)i�T�|��%�)�Wi!���7h`���4�M�Y�Åx/�.C�L]���/�*��J�ܝ1	�2j��GOV��������M����7�~��v��jҧ'Ȩ��Պn�*b�&fh�)KA6T(��Aa�ݙ�D.���o�?
�L�A�A[���S���$\s���#�֨�C���˚��T��]�kZI1�S5k]�M�F�_�ֵ&~ cMD	'���z�!Тl��@{%��o	r���ȩ�B�~<D���KZ��y�~���1���2�\��׈���e�����4���1��j�sN�#-��PN{�l�ax��Y�{�1�\�f�V��,�[0�@�ӕp C&~��4�8�j��B��)B�����-�p<�%��rz�l��Z�|Su��8����N�ZQ�m�PB>v�4skH֓�8c��>cخ壍�M�lV>pi:�����>jp�p��M�S)1�`$��$�d0��]b��	��:��8Q��L�#C�q�\�V�_ 8���	"˩�9%i'B�+�i��)F/�����T����6Z|�P���	�k<Ѵ�~j���L����
��,v��8��8~�|��?@�S�S1 _Zx�j�Y�yzU
Of�!�����+��(�#�_�o#@�5��B{���ȣJ�����;������ ����2FL������4R�� �"geͿ�#����'�!&Wi��GS�r5�)k��&@b3�`4��f��,�t� W5�5��n��#���:�����].��9�E�\�������\(���]u_K�#E�ww�Y�4�fG�G�	RK"��˲�|�O��y��(��::3��,_�.h���-��]Ü�:��4�CS1��P>�M��xB�x�x}ڎ������l
�
�x $��U��O2C��𞧿u�+��m�`��/+�`�Z�����|Z@y[�D�A��c@�̰23��e��jԾ̼�K,H�*�!N�r���Xo��D
�	O4��	1���jnt퀒��!��J����L��d�/\`8�|���a�J)���=G��b�Sl8*W���c��ćv�2{1�z�I�]U�n��_>�S&x���@ϥ�헤�� ����{ �R(�nwZ��y������^�t"���0�xY�ËG��"������$�DVnG� p��4f������ar��7�(t��]5�ct�-Yj�Ef��k%��p���)�S�������E��5g����ʏ���2���W*ϛ�@�kY���g=j�Q�{s�����p�S����(��`f74y<Ѹ*�;�t1R��L(�cx"��E���<�gUҲ�զ���fC*ѻ��9k�c6��h^]�|Zm�X�GB�ңd;s�3���ڦ}z�-�9wG���>�ڏI�o3����.�g	��(��29 �aJ�S��<���kN6騆�%��'KӴ��8�Jޢf�.fRb��|-�Di�	�bt�R-�"�~���%{ٸjRރQP���;�w=T���i����&�zK�˔-,
�ӹ�K�W˶�9�}��uV�=�m-�n=^VZ�?J5k�NM4�ϋ_0InY�w"�}li�b�eЖΈ��Xj���(bt+���8J�<u��I��h2H��Kޕ���\7�b]PPco���OO4H� ����@�ml��YO�\�\۝�Hȡ��]K`�H����$����.��8��6Kɺ��$��`�E�N(��Q�9�"؃o-g����Lh�i���� �_D�Y�5"�Y���� 1��e��Q���7�kD�C�8�F9��Q��Z�׋�Rv~�!ٳ	b6Nj��qy�qF�z"%��dF){X�/����y����oZ�{\ �0^��9>/l��Ĭ����O�+הl��=~X7�{�gO�H��t�p���!�{4�k�;�s�ݸ���el��z�n�<���U/]��}�ĸ)Ԫ�æF�8o�u.Y�I���R��\����c5������l��6�����&��6FtY�</EH_	M'��f��u}?�;%a���W*��h��Y�M֎��� ���f'm�z�����v��0N�ݧ���[sariG�����ҕ���Bl�B�%rT��PZ�TCh��/�b����G������̺� CV��3�<�n��)�%ƂU!����Ate,@����Z���!��כ���x��
p�?�)�S�[��Q�7���k�j	���	�eEJ۩�E���2ZZyd�Gw�l��AҜG0�~D��i	���|�X�*�!�_�Ӄ�Ȓq�GikU�T�^���"xȄt��,m{-}���Dab�-�Τ�h�ڡ��\�
%�%'%��0Y~����EyXh�0�wa�x�]�nvB��)�N>��Pg�؋�Z�m��{�C׶脭I�������S����3�g��D�ci9$�tM��	�Q5X�	X ��مsȲ����_^�C��4��l(ۙ����4�"ա?�g?�[��s�:�{��#���ۜ�����p�U���_!�?����̰�>s]W�$�QI�m���Pn9a�$3����B2��{Z��
�x���m��$-��ߦ�T;��� ���ī��j�ٚ"�HeJj�Ԣ��AN�Yґfl�0������C��ux+�s������})_�f�ڑ`����0�~��ہ�G|c
���rae8/�T9{i���`5V��Vg�/a ��x��j�U�|ڥ�nB��E`�Y��<=���hu�g���Z�ID��Ä�gЏ鰗�jh�$��p?Ypk:��=]��Z^,����Yw1�bY�i��nG��zT�6�Ī��r?#?D��t�<��H�
+D�J��
�J�97i1b�;��zU���������9�LLI��@f}ۤF�E}�8�*�,:=:�_�.��` ����sE�n��ې]�Sy�������_�Im<C���?�ѡ�*רʬ��(t��dK���{�:�=��س�X��5��b���Uc�SD�3mz{cu��K�j�I��9�
jZ�|���>ei�ʈ-�t��&8I�v���H�T�e\�2!>B�+��}W3(=�ΐgݾ��5�����0�F����������켉�lv�%����%������%�~�ަT\/h��Jq'��*Ҁ%o��>0�j�3���
'� (q�m�9r���}Rgf�h�Jl��>���^}?��5��`	%���GQ���k��U��AlR�v�}���ǲf��&�*Ɔ��R2�g�5�]F�V%P� ,���_뵃�C2a�<"�'ϊ��'��fur��~�]���2D����]��.T3)����v#�#�8�b��\�>s7�(�����h��&*2�d����3���TL�\��T��7ҝ1�)���6q�_6C�gŃ?[9Z��\Q�gE����U$��!T�x��H*L�thq5���!m��� �n&70��'�"�yBn<�5��0�? �vk7I�I�TL�� ��:R���M��>$�m7��3����<���u��/�M�v���1a��f}���pik���]ӎL|]�	��	�s�#S)n��XT�u�ٍ�C����!����.�$&s۪N�Q����$��;���[�!�l��������r|I3�~�zX�^4w������ 6j�r�	�i?J��[���\��y�M�Ri��h��X���?�R��U��lo��K���ܡ���'K����}��A�i�䛨���-�J�7X~�9�cD۬Roe���4'?�h�;���c}s��GD��3�����e�#\�����R_�Qh ����M�س�K/V�7o@�ըE�4� ǪV��9��w�GH��R��2��A\�T��+#�[�\��nǳ��g� 6�_��&����r>P~$�W����a�)�#^�H/�I�w=ם�� ���j-��jwHv7��b%� ?_��pb*
j����p��]
���c��*�IE�gw����\�a�?e<7:Y�,x����� ��XK3G�d��зn,Z%/�e;:��6��v���8J�hM��M�?�W�3�]Y�[���ZM��?����MC�QK=C�&�_��7Ym��c����v�.���qAol#�1�_Est�d>B�U��ȤLN#W�t���B�yV�� ��N�����O�LWl�%�gf��S"F'�^9ќ=*�0�6���
�٦��!Z_����\�b�j|.s�@�B@�f;o8_������1����B���w��d ��u����L��O��3��A�r�q�ʎj�k�>0��X��dW�yyQU�y��W���Q��G��p��
6�8.;�ٽ��3o���)�|�Q�r�B�'1��w�����˨�����5���k����ކ�l���&K4�b�O��ȗRs�z�o�=��Q�8�f��AfN45��ç<'��1�6�^��}=��|I4��1:�F�6'y���X��C��ƂCa�,-��<�7ԓ�*�՟�e��P���Ђ?3[��}?���-ό�*��u�0f��e����A�7ڽ��2z��y끕6KY�����Z�3nm���~cS�7��F˾����-1.�A!�(�Ѳ�_��boJֈ��ʹ �X�i���T���a�u]/pe�*E.�eN[n��@d�+�&���/��{W�����H�:�� �lӡ� 0i�O���g�d��� ?�/������a�jn��<��D�iu{e��R�^2Z�62�H������lv����I9cT�M�w� D�l�5v��0�+�^9���i2��/W�Q����|\)�i�+��g��*+�����v2PT��Y6�*�۰�kV�GUCI���M?��Bf#c��q�C�(,��qT�Ǿ}��J9M�S�s�����`��h���)��W�ӍI/��yk���),���//���)8=Z61b�q���ɺ�)RdK'W$��J�[�(��c��ͻ�l ��H����B���V
�9�B�r�]/��Ўc��Ty�t�u�9��^�0��y,.w��4�q�h6TR��Y�+��ڽ��)��v
�{����bTH��f��#d(ҁ_2���9�OI����FI������� � �Լ��f���-1ۈ�\{�5��k�ފ�qW[�&Z#:cnS����ϕ`~���vt1Kȸ��o�9y~�g��~U��#�w�a(l��Ѝ�]���I�%TWU����XU��ʭ����]�z��Q8�]����W�l6K�S����iv��~��m����&�_�r�u���#�r�zK='Gf�"��V��<)?1H�����������n�����CwZf`�.y׬���3�ŬȈEQ)Ep�%x���$B�7�4!���.w�3�~�w5G�P}l0nl�Ѷ�D�ë?VI��텆�v��F��cY&���j7�Um&D�j��8�X���}��S�J}��k���<�/�s�~��p'�<L�O07zʿ᜹��y��l2(��h���G2�k"FÝj�J���_�ħ�E���L"e�� ��ˑ>Ōb	��0h��[a��N�������9��I����:׈��Le(�{Z���"(C�I��C��Y-�KL�_g��v�TQ�e��";?���t �9e2q�
� �m�O���8�x��g*�����O�N?����P�G�i��_�-�?	�g �z�dRܘn����`) ��)�%�c����v�Yx0���po���D���O?p|q�CT�z�;����g?4�����K]������'o�Tl��l<��b��A���hd��qI�����g�`���|�����y`�+~C��΋��O���M��d2X���?v4�a~��$%�M�9�YUs�ڑ�x�j�ex��� {�ݯ0��EJx����YK<ԓ��h"[�A��#Y`Ltټ)�-j�f�f�Gu�5M�Y���mU�"BzW�����W���W��VQI��&�j�:�<�S��'׈��l3S���u7�S��d�5K�x�B����㥠=ǂ�O��P����̃5�R�+a ���wI���\���5�o�^~�[t^�a6r�a��Wz�*��#,:�L��� 
��<\W�k��Hu���CF�pX�;���<փ��)��MS�F�^dF_,�rg^|Ty�M鸄�Il~g��Y��4Ld�Y���~�d�0�%��.X�����BK�>d<� �����_H>P"��8]ȫAzzwO�'�Ɔ��)�]F�8d�CB��:�r��-�v��<�.d�Kc?44�����e���h�r��E�ФL�x�����ӛ�O��f3�����3����ef���*�sї�Y����*a��UQ����yd��a��r�R����fjj��'�����*j'��$,XK[}�4�I����$5�F_[?$�=�%�E(�<8�< hc�P�蒺��l<�ZU��r^!���3P��{�)*Y�h�}�~��Q�/�ln�D^�n����c48�-y�5�h���d�cZ� R�� ^{�E!aɀ�-�8��>V���|F��?�:�@.jWx��d�T̼wi��H�j����@��F�:?�����n���ie���FA1���ً� )'�5�.<�dl"&z�r�
x����g�]�n6��n��Q'�Д�Y�:�Fz���'�c�Y��3LN�6�0_ks�J�m���P	ߏ��B��\�x�j����
�|_
��;�V�&P,�T�@���ی)Fa��g����V�_�]߬	ra�i�`1 A�Dw�PRGx�g�;˿��IԠ�x�����<Yp( E�մ����C_f�Trj�6��.�m.C���F>N5ը��bC�>�-�1��"(Ӓ����:�_x3@)�(=�c�=1�gN ��y{3�8�{[������Fz@=9�:8��.Ta$UxS(v�&�˒�8�Q3��%W�.?�z�'F+7c��
��n�U���y:Y�F�Zx��f�����ے`���U�[��\�&�u�FI�΀�~��	��;���w�8��\z��/���8����w-���(�K�t���B�G�eζ���|'�.g)��Z?�����;X������+ެ�o��b����.՞l��)�y�"���>�2�����9���臾�v0|o
�*.���뾱�xL�t�	�8#07�O�mv��I�{�*<�����w���혮a��.�E:��cq׀��ZQ��9�i9n�w�n[�7nٶ�.�o`u�^��Rԗ=<�!��u:Hg쫨G|o��~>�,X��NFfyk��`� ���T��9�t�rJj�x�ά ;W*�{��*?���0���c�^�c�U�JA�9� �k�(Ô��&�����8N�B��'�B6�iL[=$ks<"{au�_?���[�M(���݅p>��ʄ�Sb�܄(���٬��+	��2�5�0�g��OHW���~��#ʽ��ę���0Dީ3<4�؀�%��,��%���'
d
��7��M�ʣ1��u��k��l����&��G�ў�@_��%WX2!RP��s�R����C���7�w�!�~0�[S�܃\����� �Ίfp�P>U�7r�^ �Mb�l���SW�8[gb飓'tI>X�P�D�i�N )��1,#��#�='�S}x�<c��0��`�7��]��Ie{���	���%���PR��"fb��6mB?�G�B��r��iʁ[�BH��3*��n{���ӷt��[zK.��݌��m���FN���w�V��w�F�-M;�+[I��!E����9�s���֎-o=n��~vk���i[� �AL�%�H��9�����(����O�A�-専	6�����A����Y�3d�ɽ"6\KH턯I��O���Dl�s<�%���5+}���HC��*�l5��?���G@=z����'Nk�TSV��T�
#C���N_�	� ���<l����K�8�������N_�8��=�N�G�*7P!���|��\��*��L��6�����81"��jA4#����xI�����Y��#}CE�Oq��>�*�r_���8�s(\��<�#b!4?�n@;ۥ�#�kK�Q:5�T�;Z�@�7��'*��
L6#���p8����x]>`OE/�֗z��	J⡡�J����L�v1<���'��Ƃ��� ��36���X_�,��jD�y�j��'�m��W��1��G@�'%z9��s��r��dBL��Q�@���Ǥ�.��U�@��w�5I���8.Bdt�{�Zv� �p���V.��6��kɆ-���Ft���.1�@朻4"ĭ�a/��>A�VeJ�f��'�e�Y���a�"��^;�'���%��f3����mH���r�v Im�R�0�̪�k�ަO�b�Ǹ]՗�w���
0g7������K�. ���!R��҃-^�kfm,X�Hhp�!�/3v6G��}��z/���)!Yl���U�a9mYq#�E��<�)�@�4U��`��L��|����n��]��=;�j�D�X���4�βP�K�����ɼ��&��20Z�1���60<) �"t��Y�D�?zg"Q�^��f�������
$��J�r�:r�g����5��K?�M"�Xo6����_��*��u}Z�w��N�
Z�V-{����x^��g�q�U��LQ���U�݁����8���L�&��`Na������Tk�J�R�E.Q��[�#�3�VP���#z��к#�8	�3��h��<k>w�ɐ]Ո�u�@�U�T��g���z�db�1|uv��V���%��>�%�sF�?���&��)��H,?����K�O�	J�������r��]�l��r��s��MkIݺR���L��;P�s�IB����ࡒ�"��$��F���<,R�Ft�ѽ`�,���0��ae��|<v旈��M}�a`�<�jCEz������S�)}6E���h&�Nf�2]H흵��3�5o�A���3���]�rٽNt��
!�NԥjK���ذ��� �·ݸ�!�r��X�8�D�تI)���l���E�#�?D�So��XGv�+K�Nl��{������ef|�������WD�P��j�j�ɷZW]L���)>Εp�V�������R9�>.���M�$9�I.�sv�7��vd���iu�����-#	�U@ke���{y˼��yB�R�"��?�c�_�jU�j|�MT��U���mAz�SXyKi֖�(<9�
�L�
�~��2��7�Ʋ8�����^\r����"�F��2�,��C�P�������ƶ��j�lx�f��Q�FqL@s�kO	���Ũ�NUf:]H��>!z��U	GG�pB�9ݿI���3\���M� �&�� �G����ԇS�G��B���z�n�u���Dz�3&�7��;W���z�)�{�F�-uQ�_i9O� G�C��gM�_%0L �a�$��j���K۰^ɾT[9���9�u<���!1�.#?�#K�=��"K�?�^���7Hͣ�7�z�-t����|�Y�����\|�}KQ�/�i�B\��jun �CD�.w�M�Qpe�.%8T'Ϻ4��)VGa��mB���p��[�e5r�588�;AJ�����b�J�s��M��0V�GWC��+E�����"����5��<�7�Z\�ɀ���v�z�e�ET�?|��y�1�a�`wO�ۙ�c̣�؏�7+��Ӊ1�$���x�4�igMI�t�U�����*46>-�ee����\��tdh>Pr<a�L�^�·��L@��8�{�����_��Kg����y5%o�^�p�Vx=��ի��n|H�o��G�_�>��)�)���^7^>&{j�
����u���0ƲW/���C
';��Jb[�o˳�^�)���� ��w��;�%v�ə0
�d4�g�h��p�~i��N ���z��HC����ad��Sm�E��Ӿl�qY�L�7�Md0�x���X��چDO�<�PE���pV�xfVN �������n$\��'��?����Ŏʛe�E��S�>���Yt����9n�:�A���ʅv�bIn���hkK�Fs�7�&�A%:膡L�e.Yߒ��W�==���h�,.$*g��#""�q�g�F>�}e���?���*�]�����c�h��"�gr28Y>d|$`~�`��J�	4����r�#5P~ͻ� eu1��ՅU�x�b@zy�жH�ؔQ��	�hPV��
�B��6-��b}M�r9(4x�##e�0����Z�.)��]���U�0�h\�	qK��}�h�?d�����>!�7\L�w z]�YF�PEB����CĴ����΃ ZyJ�l? �:�O�J�e�߆5�C�7��,e�d9*B`�q%f^����"�ҍ�}�,��g�f�5S��al�|Kؒ��kj����z�!�
�ߙ�=�vl�B�-8i��_��q����/�SG�붢��EEl��x��8��Ʒf]�I��	��t��'E�j�^�-x���0�b�� ��B�N�-��6(t�}�{ҹ�jHE�EYDڍH~Ӄ
I��j�k����2��!e ������Ft�������aG�ӂ�L`�|���`:A{cX6e���f/[��tFG�������@�'�4n�t|�5�0��B��H�W�CB���IbªH?������{uxޫK*b~?'�0��ģd��j�B�O�UA��7���,���U�+����5D"6I�g��b���X��s�������" >����^
ٷq��E��za:�c:%�ھ��Ɣ���=�R�Ԕ�my C�?ޖ��K���S,��,��1hgk]T!�>�y*�*8����fz�/Y�
�Λ%��*�,9b;�A��(���-�.8�L��vi_�� ��Si�P�W�^M�������n�X��V�d�h��?C~�;���h�f#=��a��������jbLO����`儅�8����d�N�;p ��CrO�I��"����11 o�4��,��r�Oʸ�s*�(�4	��k�y�P� �3�ė��(J#����NjL]�"=���:k�suv���YT��i��T@fd��g�T��=ȳPo�J����C�'O%O�U��̈́���^)������D��i1}�ʳ؃q{lRN?:��h�wG�?U��3(��{��;��C�b�d'R��a�
��#3�����q��_������$.�o���TUy�հ�"(��.�9�c�zvN���K�����@�|;|5�vm��r�\��so�fT3;�t��f!�b]��k{��>�zSm9	�p�D}��ç���1��nvnԽ�&�^�Ҁb*���Wƽ����/�p������(U:�T�\E�=�t�޸K�Eb	5�b�ցЙՙ���1$�GO��
������nW� �T/w�}pl���#��j��0�@G�}`�0�߽��6�� �����<⮩T�~O��a@9D�@�շ�9*��;����1�{`;1k�p^�M+7p�(&9���m�^͓9��UԹ�My��hx�r��� ��x0!4b&G�bb1K��g�(!9�dۅ�l�h|{u�xO*���;���$�d���U%�>f�ᄊ���Q��pF�#-kRQeW����	�9k�J}��^�}�{,Q�f���ճ,��T'�+�|of�S���]��X�]EA�������z�˛~l �LcGA0u�>�_� 8�*�LUo�XBt-��l���6��~V�I��$zi=�-�p8Y�&���d+�o_���]��D@էJ�u�J|hK�C�؂�〱Xo��T�\�Yꪌ�@��!��l]��=�8�����.�"���|q���6�g���%C�3��x#��_ ��ܔ�O���>���.Â�jn(��	�^Z`�f�ퟖ� ��	&��M
e1lah�0�x�ߔ�Bc.7����U�11�,�62��Rt���x�[�	ᗴ���o��a�eem�7��GLd@e^ @�`�4�rs7��;O�A�Q̬����`B�����A+_��X�CӬE��շ@H��Ɲ����ߝ�A 4��6�!O#ם&u�k��۴��{�J�LBKwS���תѲI������WW���f�������~���J4�V�8M��cSZcʸB�������5��<)0�i��]W ew:Ȩ�R平�*gf�%����[t���	?5�s1��F4`�����S?a�.�:�߱����&S�}QS����X��l6)6D�癛Jw��IR{�i����R.�E1���1E�:�TN����ͮN��h��rb.�1@@�2	��n��p��J<[�)?��i&�,��LB��[oM�7ں����~�<�y�\�T���C�'���p��DR
��=�N���Fw�x_"b��Xк�����v��5�K�M:g�D��=��P��p4�n��D���v��x�� #����@$T�����1Hl:	��%MEI@��v�jVN)���`�(��mh�<�xS�d�7��C�'ҬX�2��E�r��1w���G�2���h�~K�Pz�fRb�P��=S�0쳅��XI#��~:��Vm1�D=�!�u���{t�D�<Ƶ�C��S;���+�ц�tcMƧ�mx��x��K]G��*[p��-P������xZ�״3��K��`B����d�ﹻ��g�Sq.�������M4�jٍo�Lx^_Q4^���GV0��	)���f�>�GO*�ȇR��M�~���ܼ"��n�?�3wT
�#=Ǩ�p�'u=�c���י�~������5�fvl�-�Z��w2��2Q4Nh�KԨ~�ʐ�NV����?h���)󮙴�Ɍ ��r����q�;��$�Gg%�@���D������)�A��sU�bYS4���Z�7A��Z�ħ��l�-�W�.ڙ"E��ӝ �d��u&����{騝fIQ󾖷Ь8p}"�T`��/%��+{V�j��I�3���Ec�2~�Ic��I!r�HSӍ�\~,V$%B��H}�!�G��q���TQ�]�Ʋ��C��u�� _��Qx�T��m�yX��S�O���k�,Aߦ�����2\�a�;��Z�Y��x��Z]_��� 
�=�}q���qv.�w�u�$F8��W��!�`�-wg�1j&��:F�'��c�����q��C��7�K0p�?�����+���^�2N�he�i��F'�7ҧn����b�FHir�`�?Bқ��Ӛ���:bk_�=�����=.\������@?l�1Z�C\�
GV�聝!�X�_`U��5�;�B#S�I �y:PY~6^h�i���OP���t�uh�֕[3@GRQI�W�)����B��f�uu�5�z���9�Vqu�Om�f��$Nf��$q
��Z�������ߔaU�h���F~��a��$q��R\ ���1��ti^,�r��"�t�$΁�'������Dۢ��%��8N;E�	ņ���h��ں4e�g��X�V��7�B��~�*#��z�FS`�N_6V�D����f1�d7ca��PAA���y�o������S�./��C���ڞ���J��������TX�"���8�N�^�P�2M���.��Wji��HL�:G�#�v�g�9i>^XRDo��2Vx��BGQr���tE ��"B��'L]��Ũ���fē��M��6t��*����"����ǟv����Y�~`�X�Y陛v��x45�|x��[-.X��&����+}A�)����V��O����w4C���R!_��nO	���-�nRٙ�h��T�n����r^EԸlA�>EޒN�#?Ōb�}P�M5c���	~AU���F8ㅆ)�jK���#,T�
\��Mo.\{~!6�p�@U՝d�-�vǎ�q���D�����"�f����k��B����&�c)�v���O���������9f�ǝ8/e*A��_
� Ի�1*��:�}Z��puH;��m�����h���t!Q&f�s;�}��v�;,�[�aI!4�����Na��T��o����'v��|:�J�z"����Cv��z�Wlg���@���i���ⵗEVa� ����&^]�a�fEbo�K��HJ@u}�a�[x/'�v�K��+Ҕ�N�*���>c;��ɬ���RV�v�˔��������,�[%$l�L��@f[�I��6�_ �Stެ.%�/��9�4FQ�^��q�����2�\d�j��y �BÒ4Wc�ý�C��ݍ�`�$�k��4�W�)Gr���?��D�.�$�Z�?eP@�yb�Ź�GFE��o`V�RjG�"��k~����G�0�����L�v=�#4Y�^xwg��ɉ��~s�� �t����O�|y�j� �{	��V-����\Nd�o����;<[�,�mGr�W�D��:�=>>����͚���K8�� :�X�d�M���Rt�8���"��F��@2NvP
�qa��M�8���%����L�ipk��TS��A
���;U%��]BHi��j�2��>s�h;d��dz�������V��<��צ���$����A�*Y1�(Q�G��4`�w����2x������x���ۖ'��s���$M��9,���*m�l� �a?�� �Ora��4����g� �V�E�섐�Č;���=�I��3�}��'�DҴ~�˩�$�5DS����sUC�f ���v������ʣ>Ml߾�NSZ^&=i)lAe�̈������H��Ήح8�g�L��3������g3���h��:؇����i�+Z~L�ȸxb#���St���?�l�.�\��h:�\SG{�����o�1��Sp�.t*ʢ�?�p��aX��aNk�0�·&"Y)�}����dJ�ǜ�9�2�ߖg?�a�b�Z{n����lz����?�:�ٱq0���)�92�dB�Ԅ7�����H�l��D$L��S��}lƭ?̒4nk
�x�9b@�=�X���;��p�c��E���#�����7���'!��֥������:�5eM:bQ*�I�.��E�;�2�b[	��P*
�P+�P�k�~�0@L8^T��G�ү|�m�H"�������G�gղ�����nֺ�.�?�-�6?B�h]Vq(]��^5/�j,�n#�[�4���FL6>U��i��N��͚Vͣp����p��*����t���Tt�z��^ђx��Xg m��+����&��1QQ�*�"��5��ń�6v���b��J�$�m��Rt�����3b$�ղ�S��fF���+8'\S4���؃1��#���	�c�'��?��鿪�^��s���Yq�:��U��NV^trK�ߩ����>�\��w���M��sp��&��U���r�Rk���M��C=[V����rE�b�����ơ�>"u�v܁�����5�����K&��G�ʁ�J6�dC���i��Jb[Lpje�
s�[l/(�Y[�R����L�?��ҳ�b>Y��z�Rr��ʔ ��dל<��d$l_5��d��zz����MA���$*"d���+���NV��>	9���_z�@h4l��M��>��۔�E�Kz\�6���2��x=ß�/j�WF�7����V}D�&�Л��H|�v��\�������XP��^����h&*Z�?KP��I<�(ǈU�}�L+�u�q���Y�P]���Ap�<m�f~��������tv�H�U`>��cղ�:5�a=�8��t���q4���#��-�IH!�6�ۂ�U�l�Ď'c��J�>�= tM��<�*��'r	~�j�z��I�1�<�T�2�O�t�ϹD�?6�cC�j̮�y8��h�=nZ;My���6�td4˜��]�����-,�H"�{k����*k̺�t��u�z�ȳ���,Z�I��@q�y*#�B6��Um��'1�,zd����H����韔}�����1G�A�� ����W�w}��TU�%�C��KFس���]&i$���G0�Y`9zv9M���h!�Ge�u�h�!�5�[Bc��]� ������P�_hy��O�쭗��2o^c��a����%S�y�mؓ�7�]�i��U�J�7�����\��3�̫������5.�9��������d� ��S�,@��Zƕ-is���n4},e�Xy��|b��[	H�d�CR������r�̓�tP�V?(0���ħxjy1p�i���
�	3~�N��d��&y	�F;8e����4�Ofm.|N���� ��u�h�^��]�y@��?��6QΩ�9��^����U��K���8���H6�������F_��t�sʈ7yk�Ӱg�������P4&��R����$ r�4;�U\F^b�2�B��Q*8�ϴ���R��N	Xg�҂�vz/%i�NΪ7������,���T�ߤ?�7��#�o�eO�A�ѿX�n���)7v{p���;?,�$u "%ix� �{�>;b���Ck����R�Y��}�p�x�x��I�g�PWZ����ֆ7 ��4n�i���.u�,�T����'��F��
��?�A�htW�g#c�{R���R�
������螰W�4�h�2I��-.��';Z���^������%���˳�ۙ�e�[�����7t˙N�I���j��U`�y����������yQ`�PO'��� F� ��1{�cVt���p�\ۼ�<&�I�
�ƾ�-��F��	h�Z������|I��?'ܱe6$���7�ex���lVPlFj� S�3[���o�<q�����9���_�vuk`��J|�{3DO=o���X��g%u#H#���^?6�7��}TQc�1_-Z�"������вW^��;Ș�ck$���;��&��L	�ʆ��^Rw˰g���.\����m��g���=A٤�o���Ծ�QV7�%��㺧�e���h�V�K�|;��ƺ�G�N�&u�g�'�@5l�L�C��"K<ihG�w�p+�wk��~�ÜڂA�М��]"t�rY7�C�s\7�(c@f�C�%�H��'7������ֻ��fðzH�}�)B�E�^WE�0v�P�Y��V�Q�l��@�� fN���<6�;�oj�*�ȏ�K ����I�e}or�OysQ�5��;���5a3T�@%�L��]��[鹸k���.�Ty,�����
pg�741'���7�B� ����r0dS&�u߁»�q�(d�Pr7j3b:�hq	� �cE��+��'e�`���r��<��T��?��\�\8e�d���䕝g4�r��X����B�K&
��C�z�����?^Yܤ��z�Tq���� A'��_>�O�"j��;��w�&rv��_jɀ\���\�JX���)���!)�1tpW�qc�VwȀ�8� ����r�l���%�&�O_��ɣ�����߉�D%�X)s&kT�ZL-�S*~�>��\�}9Y$r�,6�+r�C�Pt��U
�p��QD#o!�\�`T�L�(�����>ؐFr֯W��(��BB+l}"h����,x"[�g'h�5t��	�~��&�~��*/R���x��xa$�3�x�`j�&��QBJ�M'��=Ouc����W��'�p�"�l'����d�s"�N����yX/�f�@��Z�����|��\�1���V��7L�텰��V����Î���{JpG�J��ȕIh�^'��2}&(Is�M��׹�;y���$����He�6�I��L����
�	��!'�[Sme�ЫQ�B�TҫX$�=P��+�UT���ꈢ�ۯ�,��_�6C��p_����U����@9))Cw"͞nx�7���|m�@[p�c��)^�������셶��V�ۻ��#��]�*D�ax��j��O�$�J?k�#����� �/��u#�D�x��s9�)c����#��Wx-��L�u/qQ�O�v�D�?p4Э=�
�8���]B{��?��k��H]<��zT'0=;|�ڱk���_�?ti�u�/n����3eL��Į�3��.��\�D9��yv�ZyU�)u�#g�򢠥,�FEa0��{.�1E/�nvdоh$�.���c�有ђW��s'8ą��L�{h�0+r�vAY�>:� a㠪�P����E�v(�f� �Q�_$��Rb^g땒/N�m#�+|���ڃ�_{����Rb������ұ�t��vf�����J�5�xG�g�bP��W��LJ.�����VUUT�Mv%��6�%k
�/ �!�Vh���!�?Q�`��ID\��:3K0#�`���nf)y�
��}��f/T�p��r.-�j]ˬV����W���J�{�J��u	h����T���p���8��ޣ	�?�����R^~�3e�o_.=à��)ԵL�
5-��J��ܙ��yc�"��-4��J�|��k�:"��O�bNƁ��ZqrɈ?�4#R�m�qH1�q�.󅬦������,��� �F_C_�(E���G��&TX���i���.��~�M�EI���f�A�$wA��*�:�s�Q��j��		��g����R��e�7��F��o䮑:�#��9�\ �X^�=�
cM���s�v&p� 76ޑs<�T��L����m�+�\rri�j�Y����n�,Xjv�M�Y�q&�!+O�zr"Yv��ۢ�⫞�]�pT�]�w�>č�z��F����5���.(j�O
v��ﻂQ�uY��>0kQO���6шbR�J��`[m�-%M�㚟���C����'��.)�rc"ġ�_��~��rm�[A>\8�Ȗr��7+��ʹ��}�����iL����_�lm���$#��_E��
���-&�N?8����:mIZ+��8��XqZ����z[/� �#��"��+Y�f�� `ҍ�F�h�� ��L7� �]u1����)�� ��Q�n�׃Yՙx dz;@�.�6�ݑ������@����$�Ҽ�b�j�����Z�މ����Y`�1f>AS���xmQ� �~�~�<ꛠ���}�)�I������
د�4d܌3�o���c(��u��qM}�nF�.2�TX{iL�\��:e2+���'Цfmi5��Z��P-�������X���\��po��Հ�W[���J�E�v�����~�Q ��!6U\���3x498�'oL�oF/ٟ�+J@DdL�+.�/� �*�%%�TjU�� @|�\m�Zz�N��l�o*ȁ蜽���8��Ȇ������*�'��L�2��.r��&n,x��@I�؈�R�=��ԍ����:��ԾW�7(�i���T%:��`6�kV۷ho918L�R�}C����@������?���MN��9d�Əz�#�)�R9��fi]��e��N* 	�:�/��r	�QL3/s����Z�)l~��(��{�����)�*��n�<�a�:��ocã3]��R��M��	�h�������v�����U �+��=�#�a���y¡|9����K������X�24g(�!���&����� ��p�8вE�:�����I�Z�Lȥܐ:��dм̹h�N�Dǉ��td��T|-^."Y{�PߟS�/��L����[�U��ď�p�@ލJ�BT��VJ��4��֪� ����n�;=j��F����~�ݕà��_]މ�,W���w�����68�a�!Iks� w|��n�@ݹ���"E5̀U�ɗ�ͿÉk�4
�����1�ě�U��q2��������P�.V�k$�F����$_�{m��Cf� y��!Ww>���)>a^�@�Uy	3B�d��3��ӦO޼}H�'�`��s��)_��X~Qs2C3Ř�}m��ds|n�ÊC)�?VJ��?mTx�rĢ�/-�}8poi%x�Y���y�4n<LD����urT�m4���J���90P�Q�?�����hb~��V?���R���$9z���h��Ԉb�ΖG>��΁�o����OVNNu��-R�%?�`Y�\�*7�>0�Xk���P6��Z���h8�=S���`�i\B���;�l6��.>��z���N�тܭ�ڼŬ���qWFmhZA�[IF��)��$�铃�_i@�@7�@q�C���\�]e��(�F_	P6����+�Ѷ��>���U�����a� �[qwvM$V~�ps|�^��� xZ��3 	ó�r�p����;�]FP}Խ��.���[�J��cf���q;K�0��Q��zՃ�Y���&t��ٛG�n�[z�D.�62_FZY�_�N�s:�N� �y��O��i[���y 3�\�W���: )=�@�n����M����"�뿎� ��R��O��2�hp36U+ִ�5I0e&��������<t���i�C� �O������A-�ig�ל�)D�er}%7�~�~Yf�/�
G�i�x��$����?��Ma��3m҅4�R���1B�ߠ�0��c�KH3���7�5/��0���X�L@ ʿ=s�D�9 $-{�"����RYn�s���&�CTStUD�{ř��4��`]�1����J�vjd}��:���:9�@{3�=�0N�����K�ʙtO�Q�=<!Y�A�>���XEˠ���|Y�����e�h��Λ�R` \�p�kޱvHx2�h��/W}�"F��1.[��r'q�n��A'3:g�ͳ�hś�dawrC�4�Z@��ݲ��;;c@N��zF�?�G�ք�,�Фsé��FO���d.���������*���t�*�Գʙ&*�}���'����U������B{�ga�������U���7�'��Hl}f�a܊d��y[��\�'�(7��%�ֆ]5Cu>]5��.Dde�l�w?��L���̤ `v�̖��;7�<3�*��#���	]N�<�m?�\�a��"�稔�FW
Fd� a�k\�Y��=U�[M�&���AV�Y]�y���2��K2��}����њg:\�_��q��!  ��Ɖ��;�-܂qJ��^�tє���#w�Up��4=��HR�p�B$����{"���՝�=(��,��F��s��(
�w�x��Lo�~ky�L�Ą���?��(B �LY4C�aTm�FD������yQtp�����GPk�E�3�����xgd].a�]�R�1�)��/��J�0¼��P�H�?}�O\�+���)�OP������Uxs���l���UܖE��^�>��l�z>���+l��;��P��v.� H�2��52�hrLݙNynw-�s�����I����J�}��<�1I��Q�I�يB�0���t��P�3V,����8lŋ�8t�����t�9/�K7�WD��`t��o�_N#c�UT =);�̣hQQF�(���hK`�u��vL�K���6�����S����:Eԓm�Z}U�e��aC�M"f	��&t������Q��4��Ġ��x���v���PW��ک�[p���U!?�jeGG�A��"��3CsU��G�\6 '���	M�A��JѮ�|!Ǌj���{	�'?ѿ
�_�CDa��C�KRDM8�l��m��91��#�)`yw�$�=Pئ��OU�|�
:~Dx#�KIEG5�{,��/��Y��;4���m���=B�C߮5���I?��������ۣC��5?^���uxW�(%���I�?��bp��@����%�܎�$�`^���o��I��ب���Zo�]nI�,W�Z��0^�,*_}��^��\#��>�xG��~5��s�I�n�t%ނQX�&b�czڔUP��nS��t�\�YTW�]��w�B�z���a���j%�1�c�t�V����ё���Sl�mR1#0Z���qb�.�O|�O��MO��}u'5=���7M�����3�V����,��DoE�
��I�t�.C�Y�����T�
����	=U�|V2�7��i��|�ZN����-(c4�6�g4�υ�#=5��������R����ǅ(/�?u��k���2�ꑷ0@�~��Ƽ\㺸I2�d=v�l���H�DG�r��J�9�+�H[>���ej��o�#RXX���*k=�ݯH}����J1+�V� 5�
BW���d��p�ʄ��Mc�����ê}��|/>�q�a_[��-�}sM:t�G�%�|Qy:/s�6�c�5NY;��0���$z�z4�JM��uA�,S_����q��<{hc�=���.�bw����{���9Y���-�!�$L�]���"�rФgE(2w�=�x����:9��
Y1���� ���?�#���v��1kӵ=� �r�^Z�����S�s����.+�C�u��.��w��M5��x^ڌ����5)y��Ȏ�����)��|T����3K5��͗'zV ���Ҳ�qK�/W���>�E�>�fʓ��B5���h�ac-��_��R1L�r׈���#yQ�[����Xe�٠�*&�Ix�<_T/T���i-�� gz�,g%��vB����}u�.����a���9ծ�o@Vń҉_�}�!��z�U�w�Q��7����F���.�	q}��2ea����
��ʊ�HE!q�5�;�Yp�E&�@`W�G�8՘���8�q&!0��qO9�3�FVbT7��:�r�nz+�5��Xz�]�/߫J�m���9���1��,z)�A��;qU��%�v��c�٢����ө���1�e�r�����!5�+���Lz	��ڊD��@ǈ�����O����}W=�	�˝�v�<2}��q�	�$�
X�;n�/��ך�����`D�.t<��@�!X=(�2�����n�m���R1f|b�Y��{���QP���tR�8Ė�D�χ��4!ޖ��ѝ�mh�x�K"^Q\sl�y����K�1+��ɧ��̩�U��m}�0|i�Z�F(�[�;jy���^p��Y��?mo\��f�/������3�Ã!H����v<P���;�]�T��~�b����|��R{:NT✓)�z���>˲z��>22���w7���?�)��|�Ʒ#���Oӗ�u	@�+�C�^��԰O۷d1�kX��Jba���FN�9�&;��B�c���<0�Z��Q0p���$�8V]%_~�0�6X��Y���-�;�̒�k�Sd Ü]g#'Y(�:S'�4�k����[