// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:25:51 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sN70i+rSQC95xekqi58HSXSO7CR/hJ0yOTKhQUmEUFT3IQqZVDVdVW/mhQhSzWZ7
P2+S3/549XhbLzP4TgLOgifP7sX9REZiclvBTsDwvNM8edxwcayqcSPTU6czb/A4
QSRZgkXN2bbUf/zZmf4YaFtEcr90ar0zNjmsx1AznOo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8256)
V+2LtuKl4uO4aUwtLUfZPKH2yu4VALRf/oy01qBbIBhFjkz+z0lEQWznIsfoalCx
zvlSSGPu0a4y5oTs2HIGgmxeoXY3HmfS5yPhXl1mhPFwZPUUSvBARJoPzYCRiVGd
d2hv05RkZCMwiw+I9lw7yitdXxRy0arncE9UOfbPoBiBCZRtQNrANh8peybjtg7m
b4Gp5SSwYkNljtDij0JldhYhVNKw/LzBw2ocfAbqjVZqeRHy5W1Gs18Fq2ma4o3i
10u2HYQJTCT9i0pj6iiHK53SRNJyV/0uTOWTQG6toWMIygUXth61yLl4u4vZYX66
/3LjsrJ9qmBJPfRHheNuN9njgspmohsWFSpI6vaY09Xw9vWk99lsXF4h8UlrapuS
nwPj2DEqaJhkTkUM2nNgWm+s5N8bXiQZupTKYtMjDFm/YHkr7RV1wuleJa4Ngsna
L5jPiKeixIO8DI42fnXDp/b3qwkZpLvQs+UySdaX7JNWXQKMH9z6xSZM+rId0PVX
3A9Hn3PNt4GGagpm/kDsSxNnrMqJUULsyMrqkfmNCczToulsyjnKdF/Y4j4UGpi1
aizwzqqkbaS/Xz/61yPm18e20PJtQUw4UBzyWBdkY0KmnWvjuYVorXnPAf9ArAly
Akay5QoOet5uO4XE647QtC8ewJuW0OrtD4vUhOapuEpnCMgbqxjL7XK9MRPm639P
G21KyS6rc316OHs70Yyv5q9JLjS6zZcgJ9O8y3qrEOQSd9A53rcT8lYQU8SJGGT+
sDEHsvXTcu8NR7ZPS3FI8AbVmhtOmggRcla0WSoUfpIY/NpONZtT/9X2NGCrMUMJ
KCwNZuugynJukbCiw56SOsSkP99WIQ5tKHaFdlEQdkqAt/wMzZ359MJl7NqzMLTU
4M6gpDwdSKcPs6KWrocrvqxpr18ApII5QkNTOvir4txAtUPfKwacN57J5BXQ/VbX
E8PptjkvbwV5f/YEdeq5E3xoXxlciYhmN5Xd1sj6Zv9fy0yz2oS80aThDnWnKHZm
QxHCC2Bc8qQEjprv/UbQvvMz5Mxr5ebHWCBBtDkb0wj8Gt9AuXsw95WL5J+Q6kj5
nfQ19PrSIDtDIbhRW5hsWpa7vxw4Sz8CgU+PF0kTLOZ2XEK2wjKuJ2ixMnqqnYLm
3MF/flZfxbSElJteMYIW+5JI6FjfeuQ2eql88DryOVpRkgnh1YwBeCtqZxXG6Ufw
ZSdPbgMNNGonw1j0hMnphjMJkZsqwKwlSGtsEzvp50fvQ2JvBt/YJv1TJyKSzNyZ
21A/m4orK85HnWVBM0KFJDiXbu3W6rc+a77bNlhGj0BqOtQO0EVVbsVjE5OT6Dlr
PJn3DvJ4S/s/0Nq7onggLZK4gcAe3pS6e5GC27WLZ73ercwN8GNwN/oHMb5d0AWH
hV7OLWa/14cLvQpKWUjUPrw3tIoUe+vntUWsGVSlwlsfKTMUNg2puvfh+V6JUTUL
19MSEdZG6ztICz8yYNf64g6/jYgOpdhdhsyT+AKK6MBc2b987zPv99SXP9NNUXx5
w4ysP/aoR/KlOnAERjewY1wcLSKQCw6xCO6Pvf59XbWZluKqCzbpVPA6uHChjRPn
eC1G/3a09OEgRmXdrxsEtBLNzEAbMILSjUSM1a1khqtKLtCeuSd6Y6CR/+QNzwZA
j5/qJx0+wScj2i4h4yLuiyP7horjpTAol50vrYPWR5KsOFYe1VauB0BgnHHocU/D
8n7vWcoNiwAZEwRX/WCTlXJdXp5EloRTGULEgz1Qi9CJLSWl6+WBk1EIFIVk2ySe
bGUA9AJ+vN3nbYH5c3LyLRp/d7dmKpwj8WR2C1hIls/xe0Eq8OhzWufA+L+aruOE
AbpQI8/v3Cho9kwdoaXHDU3nBaxO2mrRZMcRv0j6E/BW2RL4rfg10srpiB/1/OWC
Nqr/jBLRQKwscymufgIaY3D3n10YGCVlptpmMt7bg/TBw4BPsl+ZIf1q9774BhxV
+RL4bGhCiyT14bWIcf0bmO9gdM8CsEzFwZcT8f8jinqAaF+CZ8a7zucQTJ3uQ4wk
GwCRw9Rmh70ckDxokw+IP1Z878m1h7SZ0CDKvAUFXIwqos3qk8Fbov00mPuBdkZy
eedYfkyB4RfVWiwc1E1qHXEcVDN2ElYBOfCOW9ZV10cpM2rZTsLC6NApBEtye90L
otqYzdEisQN78yEahbsfZM70NVwIDIYf7Z1UzmwECR84dWNcITO94X+Jj9GsLxQS
FHxnTe9KQ+5fPihyqmW+hw6h9jhcWzkJcGMu9+s8gzMYeIZD/71vSQ+YgkJSWgBt
qNgeSarMa0+i/ChAPf3RUMKxr1vtjq0nwwr5MonsdAHBcQGGymRlm0avwVkArTWW
oOx0225limKXvQRS8DeDFfCn/X9hLsVXs25eqD2ye7W4pJCt2yX0mLrWwLo1r8Ha
rMc1U1+bP9H9fFzzzsYdPT/zHRv4mtUCaP6B3riKfBUNH3FNO7FJ8FxIhD3JnKpV
wcXOoFvJBCcXl+iVVPl93bvZY/mBLcsLBEFioT5rYBuDcVGI9A/eLbN11fY/4qKw
yjVNzIrdg7iJBTltemwS06/TnoV95ioGgK0/XpPcRnCIfTY8aJ3RSLExXPc/ZabR
CRLy4Fl5ytAqsmk79pditvqcTI8W1g8Hn9+uAyqkyXhQpGvJaPgtQophsZXYhU1D
VzGfX8n2SiZsrflTQFFAAK5hmMq/XCxZsQEleIIeBAWV4asy5rHIbOeYTZeAluuq
c4GVFAsIaSmEawoluMkoIH+kT1Ctw4yTykGcW62t8o8TetJrNhP6e42kTZ+SmCfj
WYi2FtYO9vgdu8rBSdBj5+fYwqQYn6pHjktaQTOm+bH4FN8bVTT41wXOZTqEnuFy
3pvYDnQWRUmc3+n1x98pP+u9buhYaC/8lZSpxODORn+8/oNSITZ+9+UPMqtsHq29
0tK/si+ZQmbRLulCume+I5KwIqNcoFIcxSnuxbUPlEao7imNfyxcTp3+cZ2Lwx/a
5gRh08cV2ErkntYdbvtIAnX8X1qSnlLbpL5lpDUqMj0gil18Rxh8NcQ0Z5mUej9i
/mgTVL6EgMgnJCud12evJg9mDdfN2jWz6edSBB77PKGiUGu6rWqyP4zjr8gNY4ES
fArXRTsQ7bDaWc6vKBMdD1Xzvf6idNAV6Z8mz5tgx370Ka9c6G5qAynQmJN/zT/o
0Ppqj2/2IxltAUjvc73p8K1hwLXtlla/OjMFA/EkAAhz1DfsWkFhM0JOdZRajl+b
PqtW6F7yylIJ28lLVhTblMl6je4LniUuMATbTsA6rg9bwz7Qzp0J6eXd1EXtRkny
66FxMS4UHHrcx857a+YkTbSUSKgCzc3ItB0Ee4+oIHWWPIZD9a0BNYZdN115itvJ
Ekzfovsr2DE2FtDjRBcnKOlJbCJHIqjF/j9zQfkdWxfrJS65UfaVUH2jj0LGsPTR
gUbLRFpiiyq7CJ4fFg81BVZVePyK0GksIGlr8QTd1a0hgJX9JB1x02rzfXQsdkYL
ym1xJ1QGK3Bzp2pVTl1MZfzODUCmpo4fR/hIGx/XM9ufrC1PVj4iqfqu0B49YGDh
2ARixSdbjp719NRhcwM8ki8n/RfN52RbV3ioZP60rcxkQr6BfkAOcgNISmK+9N1D
jfV25KkCTOzR656/Aj5jXJqU14lnWsQf9sB+vHZLGoYDYx9t2ZwnHP+rcYCC0kGV
CVgNZ1Es1OCG01SxET5cec6inKVKx3uhk6q9vF2HU5kbw/d6ohGa/ILlKDKPaCvq
1oBbtwWY+4+On6x8LLnhmM2CMxgR8bNkKKDGjxt21mO5zWHseWKA/yNTGenQJU+Z
buk9Zy6abqDuN8CUp1FdeW5nl3xU4/UesYlEMUaxZMlxoz44s4JTS2dpAeeMDF6D
JzxDDzqSqde4kYuuQw5FxFn4St/DYX01H2bhQQehB/opBvIBbSAn7R2lac/apaPA
JcfIOqBBThaGrpMEGOdXQ9vQAGgibNy0t5/pxDbfgRQL5JplaDchDIjJ66LScr0K
yi1WiR28VYT1XGZkzA8sPZE4ExLaDeTwWFNojz0M/KZ8QwweW95G2tYANvxwmKVH
TqF/BP4riSRevRHe5NeeY2x37picWbo1Xvl+w9eaMr4QT3eO7rQeAaIXNBOBzf+H
xpcANL9gRQJM4CoQT83CXKPVqTkojY9m3fd7jCqhRDIeDL0y+W59EYxg4++0GhFO
QAFbcheJuBEht3tRzkTyYV7Isphi0J4GvM+b6jENhy/j1/abrfNEoKPR8YhhOnP2
FHhMF+B9WBlB0bTBd24d6zBPt7Qz61nCdhvyXFYSGVgPK1N3PO+PryUWRWwjUY1V
cQtuhko1qdEA9sT0fW2+epnL7H7UoqBUR4d+VbothuKf/SmtPxGDKFU0uQuilUqw
C3aK24QLtaWt2PxkB34muyf6yQkXatIKPTIt8k1fH0RNKU7Flk3+flh6QOfH/FJq
TCMZ6LeIi55EZoQreeM4Sm4LHDnc9LG1VG5gFZVbOk1HfK44SjwZQGVQSrT+6Fs6
ay4bqF6pYqyndIPEt/GHOnBw4wdj7m3SXy/saC6/pv8p14kG4qII2IPdvf8D5NFC
uJS2smEhDFxQWApgS/te0OE426ZOdSpf0p16d1E6Sy1jsBGlwUoJcVyHgskESBd8
uj4hSn1tqpJACWgkpvNB5kmDasQ8oM89l0QweoC94FK1Mbbj4sqLKeeDFMUOOl3q
OwGTCRH1jxWmph9AEARzPPjXz/pXuKzqvE393l3Kvb4Uz6dWEMqAjtmfGjE+A2AK
Z43Cc2j5z6KwU9u8Q+fLZFh3AOBT0mR6mMDjBnyxnd1rJ3YONDJjy22BNPWaRlbX
wUVOG7se+Da5nstbfgrE7aWqNARS5ZnZDWJJXEuHjawIVRvOWN3jm7gRjFULLysg
HkezAAV/pdLnK3QaBkP/A6yXB7DDaaWKWOcwei3CjZwp8w610L+L8169l9YEK/2H
ZpyyTS42vqEsoSLtDUhr+Fd35sMBvCSzVAwYLaWA0iR1PeDlMmz9uje8QBW+ZKUH
qN0naFdawlnN9gl2pCMty8SuA7KWPLLaptWr0AlK5Kor6N0gk7LB1O6eT62egSsc
1wkSaaxc2d3WXRfN1xf7DgU6HuYew7lLebwrpgzPFT6J6h8EWMwgxZFKbxcitbAZ
pQ3ujJqg0ucVBkrMmum9HkyjAe47QEBRJesaXveHEIn6anTf9DXckIXdKRRSeI6v
lY6fIxroiy/nZvXzh9SHpPtL6ZcSFhMN8oTzPPem0uG5fSwz1dbBOwKuWAXvSvyf
HKj/0Ir4oHp4agXPxr8eGBcAEOzeew6tzjYwk43Vdy1oCqQ1YLR0EN6O3Bd90CgD
OgCFDLUA8aPD/EcgUfW9EO1pcPRxRILYYBZAVhidxX70xBt7oj9F4ddeo6luqvP1
x5ZyP1oQXuKjXQHCBvWs6gwCXCkP7XEXZI2VgjDEaWoVQ8ZFVxAhMspVUTZPbaBz
0MGv3eKVIMG+1pWa5F8b21+tZZla6aH3kbWP7s+ffI/oKKA+SAEagVhrWcdZqfIK
6Lm3x6wsPEXW3e6p1/otrjavDgtZkZ/r1G7KJlZMjUSIQIa/09MPTgmVPWDgfA1J
EgpUb0qrBHybkRfsg5b5jGyxsivc/TsdUvLBdi0H572rLQInJK7W/6BQJU6Hsbi7
CRbAlCh1Nj06p3iUIinYdbulz5yIJnXwi7vJLo9LDdtidn7NKPo1DRm5khobWjAX
lTI6ju74eoZRTA7msDA1d8CRR3KXxSjxF7qg0hrUa7y4HoF/EcB96kauFm9PNbSc
iiITXWh52+PbFWHSlXG/cx4hwapaNXiewX3q1wleu3BCUQ5DvBZyy6RV3xMLYFbB
rHNxqHzQBWVEbkfVtMornTyuPOMcdewgru9VPBBgmVU+fe3/fTqZkSkT7zl2JZU+
nXAdTIu8t9aMGkCs/IDh2oUKQKgNUTSVcuYCt89BiREbtUa2kL1QJd2nI6D0qGVb
rag1SixRJ7npBNtRp7ToDmj9z46n7ERr/NMCQSwZh0IOZGYvjjBA1NBIEtRmcwoP
zDEvalDJ+5onM0iNXhwP4rPYuIiNhCyTVbw9Kkl6YAecWavHWjOyzsdqwgN972d5
qfdnpPGgGfszNpPXMC/Jkk7divwjDmRgiZxbzEdIeskUxw1sEqW//kqynvLsrEll
qDUAHeWBnk3U3KOrFsKR1AYue96KdVIpDGGGQ0KPHrssKQ3jPvI+QevSyqx+7wAy
8rLQiKgA848fYqfu0USToZgZNgReAkhN+jE48I7c0/3YVI83vWlYFdTAahKtRYaI
4gtJBcplkfLApxM41PeT3Q3mwbEg7fSy1dE/Z/7wvGSEQfAKe122YV32RbF94VGu
nF9hCv2JDW5Tvaa0uJkN5NcDCdKY20pwLChO83TJBfN/+NZIX4oFXCrckntmspsp
tb5Tx8akBOwbQ0eAkvCO0Yc4tbb3tfEUeR1W5FRCuAGLG6Yn51vHHzxhqQmbtHTY
UufAc1f/Rc/dSVgx9Q68BSgChyxMaWZk8r9PhrF/+raav5VQsDBPrZ4BHxVUeSJw
/jQj+V8/8nL41uNSF/GC9u4YdID5+IAadk4RsKFl7d4503JCBSJuMR6hQWibwY4r
iwXM+e0WFv9jbOoA1sEB1OrfFfcwkWixUyDAeNcFMELYr+VsbsuG8V47qs83bG7g
y72Wq+8kKypEKxS2JLx4UFpwS4ZkeczLH4Hi4TtVT0nDnC689uXUQeUxpQVC4gIO
snw2aoeM9KI64DTNQrM9fus/PcBqh7BN37/rCXVtdV9L4XxC88i8zgI1yYomA/U2
0aDv8pE9PQtmW+6v4z6PSzNOYTGpKhKq11StHUNTFrARLS+A1Sd+hMt8legvyMsJ
Tc+ckMfgNsqUnyHt4III1IK5dc94kOb+gQACddIKMyqcUt30tqxoxjhWzclGkjwo
muKaizW+G3OHd9lVFPlsMNX7jNSqBos0b7sI9GIKyYysFI3iDZM5NsHMM8L+FLxj
Hu691J/A1wJzvtu1yWv2C/5A3HdzfJDrvFvvgKh5odChH/enRy/4xvwdaO5fZpUV
ljQ10iTKZEaElNWxsAJN6Vl6j1lpBFSjl7zgnwXL9vfgk7g/aaBkr5q1jkhsliRN
FmFWMYPVufqniQ2B8mT+rEeWQkB+JD2tbIyGtysAo+qWSgGYVihxIWmDqc5aR3BQ
qesbjh+ssa4FYzC4/qvhbeBIYCDpotBxzRD2G02g/WbdrGl1xbsNc5rvOOkELFXU
7eaYtoUe+1IrV72dQx3ZHHTkSLD+XZevdubsqbcEXYuKxqR4/cRmd0d9q1s3sEkx
R/x7V7jLpwui4RTlGcKoX59TkS8ec4Th0xOGsbsAUpHDjDHRmLJ9/a3L9ChrCBFv
eKonCQ8c2qRGd10Lq2xeezdrOutiZxtexD6vZwvul9g+SQ7u6o5h1bLO9hfA5RDB
R6VYOOGknBu5YQ3OgKHMNbMY3v/MhMbnBwUS/GsYbpdRVKyc1UIQuYejancuxjPN
xPmc6uYsg4EPK034K1XxyP9voK3h5wQcCN0Jn2y78KqRHr8h5hqsfOs2ZsXAeqse
9NBoLndfIXQvix5MjrX6nyjs6xt4jJ+vw0430wuMLzTS00VEh9T+3TmGJEwXGx3/
8DpmBN2IWINyE3I0BVM11SfxrkC1OwcQKWLEAkYnkuPvBAqMzT9fL5+nKhXLn+GL
li8cmV8fJaeZYBddXUFBDgIPbk+nAabYgN7RysFtKCvoNBUsAdhP1Cjt/dnY5EEw
X4MuCHjxAvZ4acm/r1clqxsaUYR5fPULm0n1s34eugfokPbvopXkQY+n49sHzYEN
zRoYmQp5bB7rq/+0tNHjJazmfbwLOfvWnMfSiuzruuUk4L4MWB3HQ/g5Z+d2nXO8
pcW5ndabixwvUeBw5L0gF68dzoa2geAVprvLpRJ2LcmmYWu05CtZOhHONPWihwdS
WSfp3r3GHZQTQabGYg6hkB9rflHmLLWQvhbJYFMJy93dbMPEduPI48OQkgllb2i3
J/VBIxW3xbRojVMYzPj772jAJ8jS/R4IRD8xendIpdBrzVtK5haU1ezIdZWRvRYp
0bNqdDgt+gR17Uzl8y2LFBtLBh6OzEPbGplR7gb4viRp9zPamOi9bmdoqPMZ/vL1
Qs9YHButKIzpRGTDhLbyRoDyDEwE++kebUCP97IBMGVchxzpJw8gvS3ExP5fkES1
DXBI7cJtbc93dGVkBQz/r+uR25cWMjM/Xj3E+m4ehRu6ITQmqrRH8SBBrRcBOZx9
As6U7lRRSkT74HgEqLh+D0yk3M4fAE1ha+Yr+qX6OIhEgPRNWT6iCZ8CcE3K3qje
ki0mQVylLHxveVvey4Ff3+v3jR9pEeDqoMs8LRYVH14hKKbHWZmeXv6f27lLF19d
joGhQ1X0HWrTfecr6hMAqfJtJ9TMZUn1cJ6TC4WW/FSPI2POdevxrptE80RngQus
l7FuWT0PCxF4KvKnxsgvXtLrAybu5jsjGrp1nrBVfXLsAIeV16gnALZFuUm/FM39
/KHnP7bC9+NOSGk0SxOZIzL6WFgNCG0iLhEx8enIUkJqC47t13JXL1UHO45vLrGo
zJMeCpZ8i6XIc0omdhRT4XbTAWQS9OQVDvKpKeU8qVC0xz2G0SABTBu+Vt76fRuX
yW9TLqKEdboIOQXEVoW0pLoB2LOD2/h4EClNNUFR6lgxY4wA9nJbg6FKAknO/nAY
QGaJv7Ib7Dyur2fDs3Mnw239bbp1uAHVLAfFruxTbXP55m/MHiNwIgant3UEHmVW
tP6eWyuZ8Dw7U63s5oGoMbasc0jt5l7oI1F7MRYQMRHhyoKU8HDKiQttA4TLqpL0
BDMJXTy0vUSpOBnJLX87pdXYckMfyrQzGy2kU6ZnY9PfS2Rbo3ItgO02NcA8SHPm
Y6zqeg6G4RvCa/7Wlp7YuoBMDrF4JYemNxrfouu328bQAZaJVTbwIDtiNOH3/T7F
PMeljYvhHbOKJurDBYz+MWobHD71vk8D+Xaj8XyAxw0WI79n/6jazgWECKwPOc4G
/ROBDFbdcOUQO/1cSfnZrOecUiBF3SSLz/3zaBTJX9sewxhw6SNzpMDGH0irMzMP
5Gxop0Z8n8C+thzug6KzSlis12o4gsXpKTaq1G494hO6dbPc3GP3olKk/U87QZmV
pO4I++45fbsj5seCdmMs/cbfIx6h3X0TgACF3wfrK261cDO3Rt7vzi3I42R1lg+6
s+72myEdO1T9l7sCOndPF07h1WqziCAYxKvTm1/Cg77iQPjZW8KcWmS9vn8Hvabc
uDSlIdE4jf1mD3vrkIg72uApNp08cGKKLNvfZqLYMENep0NEOgbDtrstMfATvyO+
uMZ+pPnH9+P51Fpiie2T5iQ96uNYE8ehcyV88wZekqzXupuNHTcmV/f0TEo+njIw
tgbXsDG6NUS049ZpBBXlmL40kL/r0YQtdu0LRBqfaVYTIAZu1qN6CJven0pPHzKg
wkeudasCJ/yrs4hzL7m2YUkoH7Ok9c6/9b9LGl/VgMt+BwzY3xlELtpj7AiKLB4N
oywUlV3h/cqOpNkAZns2I0eeujJzt1qyadTMwpUvDBbawAl5n79Ffki1wkE/HZ0J
CRMugV+TTVO3Ki0BLGiHtZpyqDP/8SC7jKfn2judwVxUjAJWxYMafl/CwSDm3C6o
jrea2k2YeTZsQeTlJUANc3Ct0nhV0VMa9PMMg+7aaC7mgcNV9iJFnntbYzBwbKP3
gVIkrnPjhsQbhjoHQwdOnintEC0lyB8um6auoLjCpqYYZOlIMJiDyalRXwRCbmsw
WZBHX/tVOsvBNvrafZ5DJiLn531njlHXV5CnuwRHo0vp1NyyOesMyTr4DPux25i/
5R+6RJduCifMJvOMgX1s09lrIy53nkf+j8epdpuWO7P4SO3LqmMjBU4+RC9Q5Tk+
MeUo58SSB1NIVuBEX1qwHrDq0U3rAaEk08FxEaC2zZQfrZKknhpaXgftxQhzMl7w
ckMUMgWJwYzDb/KfbSInsUioYlSR/GgjzRSpGcTqleZqCJCzU1XBg/sgeqIn7ptr
JsmbjD8qJTB7VpO5NYCW2vNppN1jzonkjf2gai0taI2xDIR3UDQ5Hbl/yuhuK0cA
WKH8jnSfRtLuF+xsBZOT9Aa4THFuAKmZDmYHRWe5wtLMNiZEluVlYnDi33oFflXG
S190392Wx2107VKF2/eA7Hh/groshbnDNV/xFSeDnYXBIWciAWTgJRyJztZzK+HB
7nAs1QQSBiS1FpekGV4lwVkdNaCd+s+i8tIV3rRLu1ZE5NQg1KQWDdTYg4VgQTu3
GkByLJ+sK7IU+iGqHaae920lQweCtDnN7yD8LSL708iURE5rDnFNtv3T1xfNzBvW
E9pSL8jxrDyIIN04y8Z+M8U4PhQgOicQkMCrGMf0uDCKhTnqX8+kHt5GYbsFPZrw
mm3vKYVRN62kJmveFeyxRfZlTsp6z/scthtS2yKEZXjy/6QHlHoQe63ZgoKmO/q1
bPM6aoxpqchaLkT9ehpaFWpAnvPg2Zue6N4jWctSm9oRMv+9Kqi6aCTMjiOMaEIa
oa1BzG09rzuCx+Hfr33ePjJURwOfiV9eqjgmfmCjNfw9WYTScQ+Uv8/TzVMn5ExW
kI1byL9oqQX4ttQtXLNXUccpBtj9B918hELFyUqpDcXq3krvRg8eSUJTFJSJz5km
IKiOnEM6LJJDueObq3PVpTcpgBCDgdPXCUnicwIbz02eElxf/jBaEFjXnlYOCiRA
AK4U6CRwtNqOsuA6XIDxZ4KWatTqYwgcV2PRHoezhttu6/1888m/jK/+yYHxx9XS
QAG8tfXrAjA86hoBGcUJswIVJcP1w50Mv5s5E7vZaxqic0xI6YkLVbpHS5rodW5r
Pmamd9o3LHtgSJAguBNjT5sFxIzJjjiKhol0Uc52llF43918n0vgOBSQA9SOg0ax
`pragma protect end_protected
